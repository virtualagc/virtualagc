// Verilog testbench created by dumbTestbench.py
`timescale 1ns / 1ps

module agc;

parameter GATE_DELAY = 20;
`include "2005267A/tb.v"

reg AGCWAR = 0, CCHG_ = 0, CDUFAL = 0, CGA17 = 0, CH1113 = 0, CH1213 = 0,
  CH1214 = 0, CH1301 = 0, CH1302 = 0, CH1303 = 0, CH1304 = 0, CH1305 = 0,
  CH1306 = 0, CH1307 = 0, CH1308 = 0, CH1309 = 0, CH1310 = 0, CH1311 = 0,
  CH1316 = 0, CH1401 = 0, CH1402 = 0, CH1403 = 0, CH1404 = 0, CH1405 = 0,
  CH1406 = 0, CH1407 = 0, CH1408 = 0, CH1409 = 0, CH1410 = 0, CH1411 = 0,
  CH1412 = 0, CH1413 = 0, CH1414 = 0, CH1416 = 0, CH3310 = 0, CH3312 = 0,
  CHWL01_ = 0, CHWL02_ = 0, CHWL03_ = 0, CHWL04_ = 0, CHWL05_ = 0, CHWL06_ = 0,
  CHWL07_ = 0, CHWL08_ = 0, CHWL09_ = 0, CHWL10_ = 0, CHWL11_ = 0, CHWL12_ = 0,
  CHWL13_ = 0, CHWL14_ = 0, CHWL16_ = 0, CTLSAT = 0, F05A_ = 0, F05B_ = 0,
  F05D = 0, FREFUN = 0, GCAPCL = 0, GOJAM = 0, GUIREL = 0, HOLFUN = 0,
  IMUCAG = 0, IMUFAL = 0, IMUOPR = 0, IN3008 = 0, IN3212 = 0, IN3213 = 0,
  IN3214 = 0, IN3216 = 0, IN3301 = 0, ISSTOR = 0, LEMATT = 0, LFTOFF = 0,
  LRRLSC = 0, LVDAGD = 0, MANRmP = 0, MANRmR = 0, MANRmY = 0, MANRpP = 0,
  MANRpR = 0, MANRpY = 0, MNIMmP = 0, MNIMmR = 0, MNIMmY = 0, MNIMpP = 0,
  MNIMpR = 0, MNIMpY = 0, OPCDFL = 0, OPMSW2 = 0, OPMSW3 = 0, OSCALM = 0,
  PCHGOF = 0, PIPAFL = 0, ROLGOF = 0, RRPONA = 0, RRRLSC = 0, S01 = 0,
  S02 = 0, S4BSAB = 0, SMSEPR = 0, SPSRDY = 0, STRPRS = 0, TEMPIN = 0,
  TPOR_ = 0, TRANmX = 0, TRANmY = 0, TRANmZ = 0, TRANpX = 0, TRANpY = 0,
  TRANpZ = 0, TRST10 = 0, TRST9 = 0, ULLTHR = 0, WCH13_ = 0, WCHG_ = 0,
  XB0_ = 0, XB1_ = 0, XB2_ = 0, XB3_ = 0, XT1_ = 0, XT3_ = 0, ZEROP = 0;

wire CCH10, CCH11, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207,
  CH3208, CH3209, CH3210, CH3313, CH3314, CH3316, CHOR01_, CHOR02_, CHOR03_,
  CHOR04_, CHOR05_, CHOR06_, CHOR07_, CHOR08_, CHOR09_, CHOR10_, CHOR11_,
  CHOR12_, CHOR13_, CHOR14_, CHOR16_, HNDRPT, RCH10_, RCH11_, RCH30_, RCH31_,
  RCH32_, RCH33_, RLYB01, RLYB02, RLYB03, RLYB04, RLYB05, RLYB06, RLYB07,
  RLYB08, RLYB09, RLYB10, RLYB11, RYWD12, RYWD13, RYWD14, RYWD16, TRP31A,
  TRP31B, TRP32, WCH10_, WCH11_, XB0;

A17 iA17 (
  rst, AGCWAR, CCHG_, CDUFAL, CGA17, CH1113, CH1213, CH1214, CH1301, CH1302,
  CH1303, CH1304, CH1305, CH1306, CH1307, CH1308, CH1309, CH1310, CH1311,
  CH1316, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406, CH1407, CH1408,
  CH1409, CH1410, CH1411, CH1412, CH1413, CH1414, CH1416, CH3310, CH3312,
  CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_, CHWL08_,
  CHWL09_, CHWL10_, CHWL11_, CHWL12_, CHWL13_, CHWL14_, CHWL16_, CTLSAT,
  F05A_, F05B_, F05D, FREFUN, GCAPCL, GOJAM, GUIREL, HOLFUN, IMUCAG, IMUFAL,
  IMUOPR, IN3008, IN3212, IN3213, IN3214, IN3216, IN3301, ISSTOR, LEMATT,
  LFTOFF, LRRLSC, LVDAGD, MANRmP, MANRmR, MANRmY, MANRpP, MANRpR, MANRpY,
  MNIMmP, MNIMmR, MNIMmY, MNIMpP, MNIMpR, MNIMpY, OPCDFL, OPMSW2, OPMSW3,
  OSCALM, PCHGOF, PIPAFL, ROLGOF, RRPONA, RRRLSC, S01, S02, S4BSAB, SMSEPR,
  SPSRDY, STRPRS, TEMPIN, TPOR_, TRANmX, TRANmY, TRANmZ, TRANpX, TRANpY,
  TRANpZ, TRST10, TRST9, ULLTHR, WCH13_, WCHG_, XB0_, XB1_, XB2_, XB3_, XT1_,
  XT3_, ZEROP, CHOR01_, CHOR02_, CHOR03_, CHOR04_, CHOR05_, CHOR06_, CHOR07_,
  CHOR08_, CHOR09_, CHOR10_, CHOR11_, CHOR12_, CHOR13_, CHOR14_, CHOR16_,
  RCH33_, XB0, CCH10, CCH11, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206,
  CH3207, CH3208, CH3209, CH3210, CH3313, CH3314, CH3316, HNDRPT, RCH10_,
  RCH11_, RCH30_, RCH31_, RCH32_, RLYB01, RLYB02, RLYB03, RLYB04, RLYB05,
  RLYB06, RLYB07, RLYB08, RLYB09, RLYB10, RLYB11, RYWD12, RYWD13, RYWD14,
  RYWD16, TRP31A, TRP31B, TRP32, WCH10_, WCH11_
);
defparam iA17.GATE_DELAY = GATE_DELAY;

endmodule
