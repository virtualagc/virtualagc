`timescale 1ns/1ps
`default_nettype none

module counter_cell_i(SIM_RST, SIM_CLK, p4VSW, GND, BKTF_n, RSSB, CA2_n, CA3_n, CA4_n, CA5_n, CXB0_n, CXB1_n, CXB2_n, CXB3_n, CXB4_n, CXB5_n, CXB6_n, CXB7_n, CG26, CDUXP, CDUXM, CDUXD, CDUYP, CDUYM, CDUYD, CDUZP, CDUZM, CDUZD, T2P, T1P, T3P, T4P, T5P, T6P, TRNP, TRNM, PIPXP, PIPXM, PIPYP, PIPYM, PIPZP, PIPZM, TRUND, SHAFTP, SHAFTM, SHAFTD, THRSTD, C32A, C32P, C32M, C33A, C33P, C33M, C24A, C25A, C26A, C34A, C34P, C34M, C35A, C35P, C35M, C27A, C30A, C31A, C40A, C40P, C40M, C41A, C41P, C41M, C53A, C54A, C55A, C36A, C36P, C36M, C37A, C37P, C37M, C50A, C51A, C52A, CG13, CG23);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire BKTF_n;
    output wire C24A;
    output wire C25A;
    output wire C26A;
    output wire C27A;
    output wire C30A;
    output wire C31A;
    output wire C32A;
    output wire C32M;
    output wire C32P;
    output wire C33A;
    output wire C33M;
    output wire C33P;
    output wire C34A;
    output wire C34M;
    output wire C34P;
    output wire C35A;
    output wire C35M;
    output wire C35P;
    output wire C36A;
    output wire C36M;
    output wire C36P;
    output wire C37A;
    output wire C37M;
    output wire C37P;
    output wire C40A;
    output wire C40M;
    output wire C40P;
    output wire C41A;
    output wire C41M;
    output wire C41P;
    output wire C50A;
    output wire C51A;
    output wire C52A;
    output wire C53A;
    output wire C54A;
    output wire C55A;
    input wire CA2_n;
    input wire CA3_n;
    input wire CA4_n;
    input wire CA5_n;
    input wire CDUXD;
    input wire CDUXM;
    input wire CDUXP;
    input wire CDUYD;
    input wire CDUYM;
    input wire CDUYP;
    input wire CDUZD;
    input wire CDUZM;
    input wire CDUZP;
    output wire CG13;
    output wire CG23;
    input wire CG26;
    input wire CXB0_n;
    input wire CXB1_n;
    input wire CXB2_n;
    input wire CXB3_n;
    input wire CXB4_n;
    input wire CXB5_n;
    input wire CXB6_n;
    input wire CXB7_n;
    input wire PIPXM;
    input wire PIPXP;
    input wire PIPYM;
    input wire PIPYP;
    input wire PIPZM;
    input wire PIPZP;
    input wire RSSB;
    input wire SHAFTD;
    input wire SHAFTM;
    input wire SHAFTP;
    input wire T1P;
    input wire T2P;
    input wire T3P;
    input wire T4P;
    input wire T5P;
    input wire T6P;
    input wire THRSTD;
    input wire TRNM;
    input wire TRNP;
    input wire TRUND;
    wire __A20_1__C10R;
    wire __A20_1__C1R;
    wire __A20_1__C2R;
    wire __A20_1__C3R;
    wire __A20_1__C4R;
    wire __A20_1__C5R;
    wire __A20_1__C6R;
    wire __A20_1__C7R;
    wire __A20_1__C8R;
    wire __A20_1__C9R;
    wire __A20_2__C10R;
    wire __A20_2__C1R;
    wire __A20_2__C2R;
    wire __A20_2__C3R;
    wire __A20_2__C4R;
    wire __A20_2__C5R;
    wire __A20_2__C6R;
    wire __A20_2__C7R;
    wire __A20_2__C8R;
    wire __A20_2__C9R;
    wire __CG11;
    wire __CG12;
    wire __CG14;
    wire __CG21;
    wire __CG22;
    wire __CG24;
    wire net_U20001_Pad1;
    wire net_U20001_Pad10;
    wire net_U20001_Pad13;
    wire net_U20001_Pad3;
    wire net_U20002_Pad10;
    wire net_U20002_Pad12;
    wire net_U20002_Pad2;
    wire net_U20002_Pad4;
    wire net_U20002_Pad5;
    wire net_U20002_Pad9;
    wire net_U20003_Pad1;
    wire net_U20003_Pad10;
    wire net_U20003_Pad13;
    wire net_U20003_Pad4;
    wire net_U20004_Pad10;
    wire net_U20004_Pad12;
    wire net_U20004_Pad13;
    wire net_U20004_Pad4;
    wire net_U20006_Pad10;
    wire net_U20006_Pad12;
    wire net_U20006_Pad13;
    wire net_U20006_Pad4;
    wire net_U20007_Pad10;
    wire net_U20007_Pad12;
    wire net_U20007_Pad13;
    wire net_U20010_Pad1;
    wire net_U20010_Pad12;
    wire net_U20010_Pad13;
    wire net_U20010_Pad3;
    wire net_U20011_Pad10;
    wire net_U20011_Pad13;
    wire net_U20011_Pad4;
    wire net_U20013_Pad1;
    wire net_U20013_Pad10;
    wire net_U20013_Pad12;
    wire net_U20013_Pad13;
    wire net_U20013_Pad3;
    wire net_U20014_Pad10;
    wire net_U20014_Pad12;
    wire net_U20014_Pad13;
    wire net_U20014_Pad4;
    wire net_U20016_Pad10;
    wire net_U20016_Pad12;
    wire net_U20016_Pad13;
    wire net_U20016_Pad4;
    wire net_U20017_Pad10;
    wire net_U20017_Pad13;
    wire net_U20019_Pad1;
    wire net_U20019_Pad10;
    wire net_U20019_Pad13;
    wire net_U20019_Pad3;
    wire net_U20020_Pad1;
    wire net_U20020_Pad10;
    wire net_U20020_Pad13;
    wire net_U20020_Pad3;
    wire net_U20022_Pad6;
    wire net_U20023_Pad3;
    wire net_U20023_Pad5;
    wire net_U20023_Pad9;
    wire net_U20024_Pad1;
    wire net_U20024_Pad10;
    wire net_U20024_Pad12;
    wire net_U20025_Pad1;
    wire net_U20025_Pad10;
    wire net_U20025_Pad12;
    wire net_U20025_Pad13;
    wire net_U20025_Pad3;
    wire net_U20026_Pad10;
    wire net_U20026_Pad12;
    wire net_U20026_Pad13;
    wire net_U20028_Pad1;
    wire net_U20028_Pad10;
    wire net_U20028_Pad13;
    wire net_U20028_Pad3;
    wire net_U20028_Pad8;
    wire net_U20030_Pad1;
    wire net_U20030_Pad10;
    wire net_U20030_Pad13;
    wire net_U20030_Pad3;
    wire net_U20031_Pad10;
    wire net_U20031_Pad12;
    wire net_U20031_Pad2;
    wire net_U20031_Pad4;
    wire net_U20031_Pad5;
    wire net_U20031_Pad9;
    wire net_U20032_Pad1;
    wire net_U20032_Pad10;
    wire net_U20032_Pad13;
    wire net_U20032_Pad4;
    wire net_U20033_Pad10;
    wire net_U20033_Pad12;
    wire net_U20033_Pad13;
    wire net_U20033_Pad4;
    wire net_U20035_Pad10;
    wire net_U20035_Pad12;
    wire net_U20035_Pad13;
    wire net_U20035_Pad4;
    wire net_U20036_Pad10;
    wire net_U20036_Pad12;
    wire net_U20036_Pad13;
    wire net_U20039_Pad1;
    wire net_U20039_Pad12;
    wire net_U20039_Pad13;
    wire net_U20039_Pad3;
    wire net_U20040_Pad10;
    wire net_U20040_Pad13;
    wire net_U20040_Pad4;
    wire net_U20042_Pad1;
    wire net_U20042_Pad10;
    wire net_U20042_Pad12;
    wire net_U20042_Pad13;
    wire net_U20042_Pad3;
    wire net_U20043_Pad10;
    wire net_U20043_Pad12;
    wire net_U20043_Pad13;
    wire net_U20043_Pad4;
    wire net_U20045_Pad10;
    wire net_U20045_Pad12;
    wire net_U20045_Pad13;
    wire net_U20045_Pad4;
    wire net_U20046_Pad10;
    wire net_U20046_Pad13;
    wire net_U20048_Pad1;
    wire net_U20048_Pad10;
    wire net_U20048_Pad13;
    wire net_U20048_Pad3;
    wire net_U20049_Pad1;
    wire net_U20049_Pad10;
    wire net_U20049_Pad13;
    wire net_U20049_Pad3;
    wire net_U20052_Pad1;
    wire net_U20052_Pad10;
    wire net_U20052_Pad12;
    wire net_U20053_Pad1;
    wire net_U20053_Pad10;
    wire net_U20053_Pad12;
    wire net_U20053_Pad13;
    wire net_U20053_Pad3;
    wire net_U20054_Pad10;
    wire net_U20054_Pad12;

    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20001(net_U20001_Pad1, CDUXP, net_U20001_Pad3, net_U20001_Pad3, net_U20001_Pad1, __A20_1__C1R, GND, CDUXM, net_U20001_Pad13, net_U20001_Pad10, net_U20001_Pad10, __A20_1__C1R, net_U20001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U20002(BKTF_n, net_U20002_Pad2, RSSB, net_U20002_Pad4, net_U20002_Pad5, __CG11, GND, __CG21, net_U20002_Pad9, net_U20002_Pad10, RSSB, net_U20002_Pad12, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20003(net_U20003_Pad1, net_U20001_Pad3, net_U20001_Pad13, net_U20003_Pad4, net_U20002_Pad2, net_U20003_Pad1, GND, net_U20003_Pad4, net_U20003_Pad13, net_U20003_Pad10, net_U20003_Pad10, __A20_1__C1R, net_U20003_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20004(C32A, __CG22, net_U20003_Pad10, net_U20004_Pad4, CDUYP, net_U20004_Pad10, GND, net_U20004_Pad4, __A20_1__C2R, net_U20004_Pad10, CDUYM, net_U20004_Pad12, net_U20004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20005(net_U20002_Pad4, CA3_n, net_U20001_Pad1, CA3_n, CXB2_n, C32P, GND, C32M, net_U20001_Pad10, CA3_n, CXB2_n, __A20_1__C1R, CXB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20006(net_U20004_Pad12, net_U20004_Pad13, __A20_1__C2R, net_U20006_Pad4, net_U20004_Pad10, net_U20004_Pad12, GND, net_U20002_Pad2, net_U20006_Pad4, net_U20006_Pad10, net_U20006_Pad10, net_U20006_Pad12, net_U20006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20007(net_U20006_Pad12, net_U20006_Pad13, __A20_1__C2R, net_U20007_Pad12, T2P, net_U20007_Pad10, GND, net_U20007_Pad12, __A20_1__C3R, net_U20007_Pad10, net_U20002_Pad2, net_U20007_Pad12, net_U20007_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20008(net_U20002_Pad4, CA3_n, net_U20004_Pad4, CA3_n, CXB3_n, C33P, GND, C33M, net_U20004_Pad13, CA3_n, CXB3_n, __A20_1__C2R, CXB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20009(__CG22, net_U20003_Pad13, __CG22, net_U20003_Pad13, net_U20006_Pad12, net_U20002_Pad5, GND, __A20_1__C3R, net_U20002_Pad4, CA2_n, CXB4_n, C33A, net_U20006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U20010(net_U20010_Pad1, net_U20007_Pad13, net_U20010_Pad3, net_U20010_Pad3, net_U20010_Pad1, __A20_1__C3R, GND, GND, net_U20010_Pad1, C24A, T1P, net_U20010_Pad12, net_U20010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20011(net_U20010_Pad12, net_U20010_Pad13, __A20_1__C4R, net_U20011_Pad4, net_U20002_Pad2, net_U20010_Pad13, GND, net_U20011_Pad4, net_U20011_Pad13, net_U20011_Pad10, net_U20011_Pad10, __A20_1__C4R, net_U20011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20012(net_U20002_Pad4, CA2_n, GND, net_U20010_Pad3, net_U20011_Pad10, C25A, GND, __A20_1__C5R, net_U20002_Pad4, CA2_n, CXB6_n, __A20_1__C4R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20013(net_U20013_Pad1, T3P, net_U20013_Pad3, net_U20013_Pad3, net_U20013_Pad1, __A20_1__C5R, GND, net_U20002_Pad2, net_U20013_Pad1, net_U20013_Pad10, net_U20013_Pad10, net_U20013_Pad12, net_U20013_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20014(net_U20013_Pad12, net_U20013_Pad13, __A20_1__C5R, net_U20014_Pad4, CDUZP, net_U20014_Pad10, GND, net_U20014_Pad4, __A20_1__C6R, net_U20014_Pad10, CDUZM, net_U20014_Pad12, net_U20014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20015(C26A, GND, net_U20010_Pad3, net_U20011_Pad13, net_U20013_Pad13,  , GND,  , GND, net_U20010_Pad3, net_U20011_Pad13, net_U20013_Pad12, net_U20002_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20016(net_U20014_Pad12, net_U20014_Pad13, __A20_1__C6R, net_U20016_Pad4, net_U20014_Pad10, net_U20014_Pad12, GND, net_U20002_Pad12, net_U20016_Pad4, net_U20016_Pad10, net_U20016_Pad10, net_U20016_Pad12, net_U20016_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20017(net_U20016_Pad12, net_U20016_Pad13, __A20_1__C6R, C34A, __CG11, net_U20016_Pad13, GND, TRNP, net_U20017_Pad13, net_U20017_Pad10, net_U20017_Pad10, __A20_1__C7R, net_U20017_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20018(net_U20002_Pad10, CA3_n, net_U20014_Pad4, CA3_n, CXB4_n, C34P, GND, C34M, net_U20014_Pad13, CA3_n, CXB4_n, __A20_1__C6R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20019(net_U20019_Pad1, TRNM, net_U20019_Pad3, net_U20019_Pad3, net_U20019_Pad1, __A20_1__C7R, GND, net_U20017_Pad13, net_U20019_Pad3, net_U20019_Pad10, net_U20002_Pad12, net_U20019_Pad10, net_U20019_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20020(net_U20020_Pad1, net_U20019_Pad13, net_U20020_Pad3, net_U20020_Pad3, net_U20020_Pad1, __A20_1__C7R, GND, T4P, net_U20020_Pad13, net_U20020_Pad10, net_U20020_Pad10, __A20_1__C8R, net_U20020_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20021(net_U20002_Pad10, CA3_n, net_U20017_Pad10, CA3_n, CXB5_n, C35P, GND, C35M, net_U20019_Pad1, CA3_n, CXB5_n, __A20_1__C7R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20022(__CG11, net_U20016_Pad12, __CG11, net_U20016_Pad12, net_U20020_Pad3, net_U20022_Pad6, GND, __A20_1__C8R, net_U20002_Pad10, CA2_n, CXB7_n, C35A, net_U20020_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U20023(net_U20022_Pad6, __CG12, net_U20023_Pad3, __CG22, net_U20023_Pad5, __CG14, GND, __CG24, net_U20023_Pad9,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20024(net_U20024_Pad1, net_U20002_Pad12, net_U20020_Pad10, net_U20024_Pad12, net_U20024_Pad1, net_U20024_Pad10, GND, net_U20024_Pad12, __A20_1__C8R, net_U20024_Pad10, __CG21, net_U20024_Pad12, C27A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20025(net_U20025_Pad1, T5P, net_U20025_Pad3, net_U20025_Pad3, net_U20025_Pad1, __A20_1__C9R, GND, net_U20002_Pad12, net_U20025_Pad1, net_U20025_Pad10, net_U20025_Pad10, net_U20025_Pad12, net_U20025_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20026(net_U20025_Pad12, net_U20025_Pad13, __A20_1__C9R, net_U20026_Pad12, T6P, net_U20026_Pad10, GND, net_U20026_Pad12, __A20_1__C10R, net_U20026_Pad10, net_U20002_Pad12, net_U20026_Pad12, net_U20026_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20027(net_U20002_Pad10, CA3_n, __CG21, net_U20024_Pad10, net_U20025_Pad13, C30A, GND, __A20_1__C10R, net_U20002_Pad10, CA3_n, CXB1_n, __A20_1__C9R, CXB0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20028(net_U20028_Pad1, net_U20026_Pad13, net_U20028_Pad3, net_U20028_Pad3, net_U20028_Pad1, __A20_1__C10R, GND, net_U20028_Pad8, net_U20028_Pad13, net_U20028_Pad10, net_U20028_Pad10, __A20_2__C10R, net_U20028_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20029(C31A, __CG21, net_U20024_Pad10, net_U20025_Pad12, net_U20028_Pad1,  , GND,  , __CG21, net_U20024_Pad10, net_U20025_Pad12, net_U20028_Pad3, net_U20023_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20030(net_U20030_Pad1, PIPYP, net_U20030_Pad3, net_U20030_Pad3, net_U20030_Pad1, __A20_2__C1R, GND, PIPYM, net_U20030_Pad13, net_U20030_Pad10, net_U20030_Pad10, __A20_2__C1R, net_U20030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U20031(BKTF_n, net_U20031_Pad2, RSSB, net_U20031_Pad4, net_U20031_Pad5, CG13, GND, CG23, net_U20031_Pad9, net_U20031_Pad10, RSSB, net_U20031_Pad12, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20032(net_U20032_Pad1, net_U20030_Pad3, net_U20030_Pad13, net_U20032_Pad4, net_U20031_Pad2, net_U20032_Pad1, GND, net_U20032_Pad4, net_U20032_Pad13, net_U20032_Pad10, net_U20032_Pad10, __A20_2__C1R, net_U20032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20033(C40A, __CG14, net_U20032_Pad10, net_U20033_Pad4, PIPZP, net_U20033_Pad10, GND, net_U20033_Pad4, __A20_2__C2R, net_U20033_Pad10, PIPZM, net_U20033_Pad12, net_U20033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20034(net_U20031_Pad4, CA4_n, net_U20030_Pad1, CA4_n, CXB0_n, C40P, GND, C40M, net_U20030_Pad10, CA4_n, CXB0_n, __A20_2__C1R, CXB0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20035(net_U20033_Pad12, net_U20033_Pad13, __A20_2__C2R, net_U20035_Pad4, net_U20033_Pad10, net_U20033_Pad12, GND, net_U20031_Pad2, net_U20035_Pad4, net_U20035_Pad10, net_U20035_Pad10, net_U20035_Pad12, net_U20035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20036(net_U20035_Pad12, net_U20035_Pad13, __A20_2__C2R, net_U20036_Pad12, TRUND, net_U20036_Pad10, GND, net_U20036_Pad12, __A20_2__C3R, net_U20036_Pad10, net_U20031_Pad2, net_U20036_Pad12, net_U20036_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20037(net_U20031_Pad4, CA4_n, net_U20033_Pad4, CA4_n, CXB1_n, C41P, GND, C41M, net_U20033_Pad13, CA4_n, CXB1_n, __A20_2__C2R, CXB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20038(__CG14, net_U20032_Pad13, __CG14, net_U20032_Pad13, net_U20035_Pad12, net_U20031_Pad5, GND, __A20_2__C3R, net_U20031_Pad4, CA5_n, CXB3_n, C41A, net_U20035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U20039(net_U20039_Pad1, net_U20036_Pad13, net_U20039_Pad3, net_U20039_Pad3, net_U20039_Pad1, __A20_2__C3R, GND, __CG24, net_U20039_Pad1, C53A, SHAFTD, net_U20039_Pad12, net_U20039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20040(net_U20039_Pad12, net_U20039_Pad13, __A20_2__C4R, net_U20040_Pad4, net_U20031_Pad2, net_U20039_Pad13, GND, net_U20040_Pad4, net_U20040_Pad13, net_U20040_Pad10, net_U20040_Pad10, __A20_2__C4R, net_U20040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20041(net_U20031_Pad4, CA5_n, __CG24, net_U20039_Pad3, net_U20040_Pad10, C54A, GND, __A20_2__C5R, net_U20031_Pad4, CA5_n, CXB5_n, __A20_2__C4R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20042(net_U20042_Pad1, THRSTD, net_U20042_Pad3, net_U20042_Pad3, net_U20042_Pad1, __A20_2__C5R, GND, net_U20031_Pad2, net_U20042_Pad1, net_U20042_Pad10, net_U20042_Pad10, net_U20042_Pad12, net_U20042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20043(net_U20042_Pad12, net_U20042_Pad13, __A20_2__C5R, net_U20043_Pad4, SHAFTP, net_U20043_Pad10, GND, net_U20043_Pad4, __A20_2__C6R, net_U20043_Pad10, SHAFTM, net_U20043_Pad12, net_U20043_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20044(C55A, __CG24, net_U20039_Pad3, net_U20040_Pad13, net_U20042_Pad13,  , GND,  , __CG24, net_U20039_Pad3, net_U20040_Pad13, net_U20042_Pad12, net_U20031_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20045(net_U20043_Pad12, net_U20043_Pad13, __A20_2__C6R, net_U20045_Pad4, net_U20043_Pad10, net_U20043_Pad12, GND, net_U20031_Pad12, net_U20045_Pad4, net_U20045_Pad10, net_U20045_Pad10, net_U20045_Pad12, net_U20045_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20046(net_U20045_Pad12, net_U20045_Pad13, __A20_2__C6R, C36A, __CG12, net_U20045_Pad13, GND, PIPXP, net_U20046_Pad13, net_U20046_Pad10, net_U20046_Pad10, __A20_2__C7R, net_U20046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20047(net_U20031_Pad10, CA3_n, net_U20043_Pad4, CA3_n, CXB6_n, C36P, GND, C36M, net_U20043_Pad13, CA3_n, CXB6_n, __A20_2__C6R, CXB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20048(net_U20048_Pad1, PIPXM, net_U20048_Pad3, net_U20048_Pad3, net_U20048_Pad1, __A20_2__C7R, GND, net_U20046_Pad13, net_U20048_Pad3, net_U20048_Pad10, net_U20031_Pad12, net_U20048_Pad10, net_U20048_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20049(net_U20049_Pad1, net_U20048_Pad13, net_U20049_Pad3, net_U20049_Pad3, net_U20049_Pad1, __A20_2__C7R, GND, CDUXD, net_U20049_Pad13, net_U20049_Pad10, net_U20049_Pad10, __A20_2__C8R, net_U20049_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20050(net_U20031_Pad10, CA3_n, net_U20046_Pad10, CA3_n, CXB7_n, C37P, GND, C37M, net_U20048_Pad1, CA3_n, CXB7_n, __A20_2__C7R, CXB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20051(__CG12, net_U20045_Pad12, __CG12, net_U20045_Pad12, net_U20049_Pad3, net_U20023_Pad5, GND, __A20_2__C8R, net_U20031_Pad10, CA5_n, CXB0_n, C37A, net_U20049_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20052(net_U20052_Pad1, net_U20031_Pad12, net_U20049_Pad10, net_U20052_Pad12, net_U20052_Pad1, net_U20052_Pad10, GND, net_U20052_Pad12, __A20_2__C8R, net_U20052_Pad10, CG26, net_U20052_Pad12, C50A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20053(net_U20053_Pad1, CDUYD, net_U20053_Pad3, net_U20053_Pad3, net_U20053_Pad1, __A20_2__C9R, GND, net_U20031_Pad12, net_U20053_Pad1, net_U20053_Pad10, net_U20053_Pad10, net_U20053_Pad12, net_U20053_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20054(net_U20053_Pad12, net_U20053_Pad13, __A20_2__C9R, net_U20054_Pad12, CDUZD, net_U20054_Pad10, GND, net_U20054_Pad12, __A20_2__C10R, net_U20054_Pad10, net_U20031_Pad12, net_U20054_Pad12, net_U20028_Pad8, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20055(net_U20031_Pad10, CA5_n, CG26, net_U20052_Pad10, net_U20053_Pad13, C51A, GND, __A20_2__C10R, net_U20031_Pad10, CA5_n, CXB2_n, __A20_2__C9R, CXB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20056(C52A, CG26, net_U20052_Pad10, net_U20053_Pad12, net_U20028_Pad10,  , GND,  , CG26, net_U20052_Pad10, net_U20053_Pad12, net_U20028_Pad13, net_U20023_Pad9, p4VSW, SIM_RST, SIM_CLK);
endmodule