// Verilog testbench created by dumbTestbench.py
`timescale 100ns / 1ns

module agc;

reg rst = 1;
reg STRT2 = 1;
initial
  begin
    $dumpfile("agc.lxt2");
    $dumpvars(0, agc);
    # 1 rst = 0;
    # 50 STRT2 = 0;
    # 1000 $finish;
  end

reg CLOCK = 0;
always #2.44140625 CLOCK = !CLOCK;

reg BR1B2B = 0, BR2_ = 0, CGA3 = 0, CT_ = 0, DBLTST = 0, EXT = 0, EXTPLS = 0,
  FS09 = 0, FS10 = 0, GOJAM = 0, INHPLS = 0, INKL = 0, KRPT = 0, MNHRPT = 0,
  MTCSAI = 0, NISQ = 0, ODDSET_ = 0, OVNHRP = 0, PHS2_ = 0, RELPLS = 0,
  RT_ = 0, RUPTOR_ = 0, RXOR0 = 0, ST0_ = 0, ST1_ = 0, ST3_ = 0, STD2 = 0,
  T01_ = 0, T02 = 0, T07DC_ = 0, T12_ = 0, WL10_ = 0, WL11_ = 0, WL12_ = 0,
  WL13_ = 0, WL14_ = 0, WL16_ = 0, WT_ = 0, d5XP4 = 0;

wire AD0, ADS0, AUG0, AUG0_, BMF0, BMF0_, BZF0, BZF0_, CCS0, CCS0_, CON1,
  CON2, CSQG, DAS0, DAS0_, DAS1, DAS1_, DCA0, DCS0, DIM0, DIM0_, DXCH0,
  EXST0_, EXST1_, FUTEXT, GOJ1, GOJ1_, IC1, IC10, IC10_, IC11, IC12, IC12_,
  IC13, IC13_, IC14, IC15, IC15_, IC16, IC16_, IC17, IC2, IC2_, IC3, IC3_,
  IC4, IC4_, IC5, IC5_, IC6, IC7, IC8_, IC9, IC9_, IIP, IIP_, INCR0, INHINT,
  INKBT1, LXCH0, MASK0, MASK0_, MIIP, MINHL, MP0, MP0_, MP1, MP1_, MP3,
  MP3_, MSQ10, MSQ11, MSQ12, MSQ13, MSQ14, MSQ16, MSQEXT, MSU0, MSU0_,
  MTCSA_, NDX0, NDX0_, NDXX1, NDXX1_, NEXST0, NEXST0_, NISQL_, QC0, QC0_,
  QC1_, QC2_, QC3_, QXCH0, QXCH0_, RBSQ, RPTFRC, RPTSET, RSM3, RSM3_, SCAS10,
  SQ0_, SQ1_, SQ2_, SQ3_, SQ4_, SQ5, SQ5QC0_, SQ5_, SQ6_, SQ7_, SQEXT,
  SQEXT_, SQR10, SQR10_, SQR11, SQR12, SQR12_, SQR13, SQR14, SQR16, STRTFC,
  SU0, T07, TC0, TC0_, TCF0, TCSAJ3, TCSAJ3_, TS0, TS0_, WSQG_;

A3 iA3 (
  rst, BR1B2B, BR2_, CGA3, CT_, DBLTST, EXT, EXTPLS, FS09, FS10, GOJAM, INHPLS,
  INKL, KRPT, MNHRPT, MTCSAI, NISQ, ODDSET_, OVNHRP, PHS2_, RELPLS, RT_,
  RUPTOR_, RXOR0, ST0_, ST1_, ST3_, STD2, T01_, T02, T07DC_, T12_, WL10_,
  WL11_, WL12_, WL13_, WL14_, WL16_, WT_, d5XP4, CON1, CON2, EXST0_, INKBT1,
  MIIP, MINHL, MSQ10, MSQ11, MSQ12, MSQ13, MSQ14, MSQ16, MSQEXT, MTCSA_,
  NEXST0, QC0, QC0_, QC1_, QC2_, QC3_, RPTSET, SCAS10, SQ0_, SQ1_, SQ2_,
  SQ3_, SQ4_, SQ5, SQ6_, SQ7_, SQEXT, SQEXT_, T07, TCSAJ3, TS0, AD0, ADS0,
  AUG0, AUG0_, BMF0, BMF0_, BZF0, BZF0_, CCS0, CCS0_, CSQG, DAS0, DAS0_,
  DAS1, DAS1_, DCA0, DCS0, DIM0, DIM0_, DXCH0, EXST1_, FUTEXT, GOJ1, GOJ1_,
  IC1, IC10, IC10_, IC11, IC12, IC12_, IC13, IC13_, IC14, IC15, IC15_, IC16,
  IC16_, IC17, IC2, IC2_, IC3, IC3_, IC4, IC4_, IC5, IC5_, IC6, IC7, IC8_,
  IC9, IC9_, IIP, IIP_, INCR0, INHINT, LXCH0, MASK0, MASK0_, MP0, MP0_, MP1,
  MP1_, MP3, MP3_, MSU0, MSU0_, NDX0, NDX0_, NDXX1, NDXX1_, NEXST0_, NISQL_,
  QXCH0, QXCH0_, RBSQ, RPTFRC, RSM3, RSM3_, SQ5QC0_, SQ5_, SQR10, SQR10_,
  SQR11, SQR12, SQR12_, SQR13, SQR14, SQR16, STRTFC, SU0, TC0, TC0_, TCF0,
  TCSAJ3_, TS0_, WSQG_
);

initial $timeformat(-9, 0, " ns", 10);
initial $monitor("%t: %d", $time, CLOCK);

endmodule
