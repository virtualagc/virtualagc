`timescale 1ns/1ps
`default_nettype none

module four_bit_2(SIM_RST, SIM_CLK, p4VSW, GND, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI05_n, CO06, MONEX, XUY09_n, XUY10_n, CH05, CH06, CH07, CH08, G05ED, G06ED, G07ED, L04_n, G2LSG_n, G09_n, G10_n, G11_n, MDT05, MDT06, MDT07, MDT08, SA05, SA06, SA07, SA08, RBLG_n, RULOG_n, WL09_n, WL10_n, WG1G_n, WG3G_n, WG4G_n, WYDG_n, WYLOG_n, R1C, WL04_n, WHOMP, CI09_n, CO10, G05, G05_n, G06, G06_n, G07, G07_n, G08, L08_n, RL05_n, RL06_n, XUY05_n, XUY06_n, WL05, WL05_n, WL06, WL06_n, WL07, WL07_n, WL08, WL08_n, GEM05, GEM06, GEM07, GEM08, MWL05, MWL06, MWL07, MWL08);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire A2XG_n;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH05;
    input wire CH06;
    input wire CH07;
    input wire CH08;
    input wire CI05_n;
    output wire CI09_n;
    input wire CLG1G;
    input wire CLXC;
    input wire CO06;
    output wire CO10; //FPGA#wand
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire G05;
    input wire G05ED;
    inout wire G05_n; //FPGA#wand
    output wire G06;
    input wire G06ED;
    inout wire G06_n; //FPGA#wand
    output wire G07;
    input wire G07ED;
    inout wire G07_n; //FPGA#wand
    output wire G08;
    input wire G09_n;
    input wire G10_n;
    input wire G11_n;
    input wire G2LSG_n;
    output wire GEM05;
    output wire GEM06;
    output wire GEM07;
    output wire GEM08;
    input wire L04_n;
    inout wire L08_n; //FPGA#wand
    input wire L2GDG_n;
    input wire MDT05;
    input wire MDT06;
    input wire MDT07;
    input wire MDT08;
    input wire MONEX;
    output wire MWL05; //FPGA#wand
    output wire MWL06; //FPGA#wand
    output wire MWL07; //FPGA#wand
    output wire MWL08; //FPGA#wand
    input wire R1C;
    input wire RAG_n;
    input wire RBLG_n;
    input wire RCG_n;
    input wire RGG_n;
    inout wire RL05_n; //FPGA#wand
    inout wire RL06_n; //FPGA#wand
    input wire RLG_n;
    input wire RQG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA05;
    input wire SA06;
    input wire SA07;
    input wire SA08;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WHOMP;
    input wire WL04_n;
    output wire WL05;
    output wire WL05_n;
    output wire WL06;
    output wire WL06_n;
    output wire WL07;
    output wire WL07_n;
    output wire WL08;
    output wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYLOG_n;
    input wire WZG_n;
    output wire XUY05_n;
    output wire XUY06_n;
    input wire XUY09_n;
    input wire XUY10_n;
    wire __A09_1__X1;
    wire __A09_1__X1_n;
    wire __A09_1__X2;
    wire __A09_1__X2_n;
    wire __A09_1__Y1;
    wire __A09_1__Y1_n;
    wire __A09_1__Y2;
    wire __A09_1__Y2_n;
    wire __A09_1___A1_n;
    wire __A09_1___A2_n;
    wire __A09_1___B1_n;
    wire __A09_1___B2_n;
    wire __A09_1___CI_INTERNAL;
    wire __A09_1___Q1_n;
    wire __A09_1___Q2_n;
    wire __A09_1___RL_OUT_1;
    wire __A09_1___RL_OUT_2;
    wire __A09_1___SUMA1;
    wire __A09_1___SUMA2;
    wire __A09_1___SUMB1;
    wire __A09_1___SUMB2;
    wire __A09_1___Z1_n; //FPGA#wand
    wire __A09_1___Z2_n; //FPGA#wand
    wire __A09_2__X1;
    wire __A09_2__X1_n;
    wire __A09_2__X2;
    wire __A09_2__X2_n;
    wire __A09_2__Y1;
    wire __A09_2__Y1_n;
    wire __A09_2__Y2;
    wire __A09_2__Y2_n;
    wire __A09_2___A1_n;
    wire __A09_2___A2_n;
    wire __A09_2___B1_n;
    wire __A09_2___B2_n;
    wire __A09_2___CI_INTERNAL;
    wire __A09_2___Q1_n;
    wire __A09_2___Q2_n;
    wire __A09_2___RL1_n; //FPGA#wand
    wire __A09_2___RL2_n; //FPGA#wand
    wire __A09_2___RL_OUT_1;
    wire __A09_2___RL_OUT_2;
    wire __A09_2___SUMA1;
    wire __A09_2___SUMA2;
    wire __A09_2___SUMB1;
    wire __A09_2___SUMB2;
    wire __A09_2___Z1_n; //FPGA#wand
    wire __A09_2___Z2_n; //FPGA#wand
    wire __CI07_n;
    wire __CO08; //FPGA#wand
    wire __G08_n; //FPGA#wand
    wire __L05_n; //FPGA#wand
    wire __L06_n; //FPGA#wand
    wire __L07_n; //FPGA#wand
    wire __XUY07_n;
    wire __XUY08_n;
    wire net_U9001_Pad1;
    wire net_U9001_Pad10;
    wire net_U9001_Pad4;
    wire net_U9003_Pad1;
    wire net_U9003_Pad10;
    wire net_U9004_Pad1;
    wire net_U9004_Pad12;
    wire net_U9004_Pad13;
    wire net_U9004_Pad2;
    wire net_U9004_Pad6;
    wire net_U9004_Pad8;
    wire net_U9005_Pad12;
    wire net_U9005_Pad2;
    wire net_U9006_Pad10;
    wire net_U9006_Pad13;
    wire net_U9006_Pad4;
    wire net_U9007_Pad11;
    wire net_U9007_Pad13;
    wire net_U9007_Pad3;
    wire net_U9007_Pad5;
    wire net_U9007_Pad9;
    wire net_U9008_Pad1;
    wire net_U9008_Pad10;
    wire net_U9008_Pad13;
    wire net_U9008_Pad4;
    wire net_U9009_Pad1;
    wire net_U9009_Pad13;
    wire net_U9009_Pad4;
    wire net_U9010_Pad1;
    wire net_U9010_Pad13;
    wire net_U9010_Pad4;
    wire net_U9011_Pad10;
    wire net_U9011_Pad11;
    wire net_U9011_Pad13;
    wire net_U9011_Pad8;
    wire net_U9011_Pad9;
    wire net_U9012_Pad13;
    wire net_U9012_Pad4;
    wire net_U9013_Pad1;
    wire net_U9013_Pad11;
    wire net_U9013_Pad13;
    wire net_U9013_Pad5;
    wire net_U9013_Pad9;
    wire net_U9014_Pad10;
    wire net_U9014_Pad13;
    wire net_U9016_Pad1;
    wire net_U9016_Pad4;
    wire net_U9018_Pad11;
    wire net_U9018_Pad12;
    wire net_U9018_Pad13;
    wire net_U9019_Pad1;
    wire net_U9019_Pad10;
    wire net_U9019_Pad4;
    wire net_U9021_Pad1;
    wire net_U9021_Pad13;
    wire net_U9022_Pad1;
    wire net_U9022_Pad12;
    wire net_U9022_Pad8;
    wire net_U9023_Pad10;
    wire net_U9023_Pad13;
    wire net_U9023_Pad4;
    wire net_U9024_Pad10;
    wire net_U9024_Pad11;
    wire net_U9024_Pad4;
    wire net_U9024_Pad9;
    wire net_U9026_Pad4;
    wire net_U9026_Pad5;
    wire net_U9026_Pad6;
    wire net_U9026_Pad8;
    wire net_U9027_Pad1;
    wire net_U9027_Pad10;
    wire net_U9028_Pad13;
    wire net_U9028_Pad3;
    wire net_U9028_Pad9;
    wire net_U9029_Pad1;
    wire net_U9029_Pad10;
    wire net_U9030_Pad1;
    wire net_U9030_Pad10;
    wire net_U9030_Pad13;
    wire net_U9031_Pad13;
    wire net_U9031_Pad2;
    wire net_U9031_Pad3;
    wire net_U9031_Pad4;
    wire net_U9031_Pad8;
    wire net_U9035_Pad1;
    wire net_U9035_Pad10;
    wire net_U9035_Pad4;
    wire net_U9037_Pad1;
    wire net_U9037_Pad10;
    wire net_U9038_Pad1;
    wire net_U9038_Pad12;
    wire net_U9038_Pad2;
    wire net_U9038_Pad6;
    wire net_U9038_Pad8;
    wire net_U9039_Pad12;
    wire net_U9039_Pad2;
    wire net_U9040_Pad10;
    wire net_U9040_Pad13;
    wire net_U9040_Pad4;
    wire net_U9041_Pad11;
    wire net_U9041_Pad13;
    wire net_U9041_Pad3;
    wire net_U9041_Pad5;
    wire net_U9041_Pad9;
    wire net_U9042_Pad10;
    wire net_U9042_Pad11;
    wire net_U9042_Pad4;
    wire net_U9042_Pad9;
    wire net_U9044_Pad1;
    wire net_U9044_Pad6;
    wire net_U9045_Pad13;
    wire net_U9045_Pad4;
    wire net_U9046_Pad1;
    wire net_U9046_Pad13;
    wire net_U9046_Pad4;
    wire net_U9047_Pad1;
    wire net_U9047_Pad13;
    wire net_U9047_Pad4;
    wire net_U9048_Pad1;
    wire net_U9048_Pad10;
    wire net_U9048_Pad13;
    wire net_U9048_Pad4;
    wire net_U9049_Pad11;
    wire net_U9049_Pad8;
    wire net_U9050_Pad11;
    wire net_U9050_Pad13;
    wire net_U9050_Pad5;
    wire net_U9052_Pad11;
    wire net_U9052_Pad12;
    wire net_U9052_Pad13;
    wire net_U9053_Pad1;
    wire net_U9053_Pad10;
    wire net_U9053_Pad4;
    wire net_U9055_Pad13;
    wire net_U9056_Pad10;
    wire net_U9056_Pad13;
    wire net_U9056_Pad4;
    wire net_U9057_Pad10;
    wire net_U9057_Pad11;
    wire net_U9057_Pad4;
    wire net_U9057_Pad9;
    wire net_U9059_Pad4;
    wire net_U9059_Pad5;
    wire net_U9059_Pad6;
    wire net_U9059_Pad8;
    wire net_U9060_Pad1;
    wire net_U9060_Pad10;
    wire net_U9061_Pad3;
    wire net_U9062_Pad1;
    wire net_U9062_Pad10;
    wire net_U9063_Pad1;
    wire net_U9063_Pad10;

    pullup R9001(__CO08);
    pullup R9002(RL05_n);
    pullup R9003(__L05_n);
    pullup R9005(__A09_1___Z1_n);
    pullup R9006(G05_n);
    pullup R9007(RL06_n);
    pullup R9008(__L06_n);
    pullup R9009(__A09_1___Z2_n);
    pullup R9010(G06_n);
    pullup R9011(CO10);
    pullup R9012(__A09_2___RL1_n);
    pullup R9013(__L07_n);
    pullup R9015(__A09_2___Z1_n);
    pullup R9016(G07_n);
    pullup R9017(__A09_2___RL2_n);
    pullup R9018(L08_n);
    pullup R9019(__A09_2___Z2_n);
    pullup R9020(__G08_n);
    U74HC02 U9001(net_U9001_Pad1, A2XG_n, __A09_1___A1_n, net_U9001_Pad4, WYLOG_n, WL05_n, GND, WL04_n, WYDG_n, net_U9001_Pad10, __A09_1__Y1_n, CUG, __A09_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9002(MONEX, net_U9001_Pad1, __A09_1__X1_n, CLXC, CUG, __A09_1__X1, GND, __A09_1__Y1_n, net_U9001_Pad4, net_U9001_Pad10, __A09_1__Y1, __A09_1__X1_n, __A09_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9003(net_U9003_Pad1, __A09_1__X1_n, __A09_1__Y1_n, XUY05_n, __A09_1__X1, __A09_1__Y1, GND, net_U9003_Pad1, XUY05_n, net_U9003_Pad10, net_U9003_Pad1, __A09_1___SUMA1, __A09_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9004(net_U9004_Pad1, net_U9004_Pad2, __A09_1___SUMA1, __A09_1___SUMB1, RULOG_n, net_U9004_Pad6, GND, net_U9004_Pad8, __XUY07_n, XUY05_n, CI05_n, net_U9004_Pad12, net_U9004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9005(CI05_n, net_U9005_Pad2, G05_n, GEM05, RL05_n, WL05, GND, WL05_n, WL05,  ,  , net_U9005_Pad12, __A09_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9006(__A09_1___SUMB1, net_U9003_Pad10, net_U9005_Pad2, net_U9006_Pad4, WAG_n, WL05_n, GND, WL07_n, WALSG_n, net_U9006_Pad10, __A09_1___A1_n, CAG, net_U9006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9007(net_U9004_Pad8, __CO08, net_U9007_Pad3, RL05_n, net_U9007_Pad5, __L05_n, GND, __A09_1___Z1_n, net_U9007_Pad9, RL05_n, net_U9007_Pad11, RL05_n, net_U9007_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U9008(net_U9008_Pad1, RAG_n, __A09_1___A1_n, net_U9008_Pad4, WLG_n, WL05_n, GND, __G08_n, G2LSG_n, net_U9008_Pad10, __L05_n, CLG1G, net_U9008_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9009(net_U9009_Pad1, WG1G_n, WL08_n, net_U9009_Pad4, WQG_n, WL05_n, GND, net_U9009_Pad4, net_U9009_Pad13, __A09_1___Q1_n, __A09_1___Q1_n, CQG, net_U9009_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9010(net_U9010_Pad1, RQG_n, __A09_1___Q1_n, net_U9010_Pad4, WZG_n, WL05_n, GND, net_U9010_Pad4, net_U9010_Pad13, net_U9007_Pad9, __A09_1___Z1_n, CZG, net_U9010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9011(__A09_1___RL_OUT_1, net_U9010_Pad1, MDT05, R1C, GND, net_U9007_Pad13, GND, net_U9011_Pad8, net_U9011_Pad9, net_U9011_Pad10, net_U9011_Pad11, net_U9007_Pad11, net_U9011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9012(net_U9011_Pad13, RZG_n, __A09_1___Z1_n, net_U9012_Pad4, WBG_n, WL05_n, GND, net_U9012_Pad4, net_U9012_Pad13, __A09_1___B1_n, __A09_1___B1_n, CBG, net_U9012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9013(net_U9013_Pad1, __CO08, net_U9011_Pad8, RL05_n, net_U9013_Pad5, G05_n, GND, G05_n, net_U9013_Pad9, RL06_n, net_U9013_Pad11, __L06_n, net_U9013_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U9014(net_U9011_Pad9, RBLG_n, __A09_1___B1_n, net_U9011_Pad10, net_U9012_Pad13, RCG_n, GND, WL04_n, WG3G_n, net_U9014_Pad10, WL06_n, WG4G_n, net_U9014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9015(net_U9006_Pad4, net_U9006_Pad10, net_U9004_Pad6, net_U9008_Pad1, CH05, net_U9007_Pad3, GND, net_U9007_Pad5, net_U9008_Pad4, net_U9008_Pad10, net_U9008_Pad13, __A09_1___A1_n, net_U9006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9016(net_U9016_Pad1, L2GDG_n, L04_n, net_U9016_Pad4, WG1G_n, WL05_n, GND, G05_n, CGG, G05, RGG_n, G05_n, net_U9011_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9017(net_U9016_Pad1, net_U9016_Pad4, GND, __XUY08_n, XUY06_n, net_U9013_Pad1, GND, __A09_1___RL_OUT_1, RLG_n, __L05_n, GND, net_U9013_Pad9, G05, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U9018(net_U9013_Pad5, G05ED, SA05, net_U9014_Pad10, net_U9014_Pad13,  , GND,  , G06ED, SA06, net_U9018_Pad11, net_U9018_Pad12, net_U9018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9019(net_U9019_Pad1, A2XG_n, __A09_1___A2_n, net_U9019_Pad4, WYLOG_n, WL06_n, GND, WL05_n, WYDG_n, net_U9019_Pad10, __A09_1__Y2_n, CUG, __A09_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9020(MONEX, net_U9019_Pad1, __A09_1__X2_n, CLXC, CUG, __A09_1__X2, GND, __A09_1__Y2_n, net_U9019_Pad4, net_U9019_Pad10, __A09_1__Y2, __A09_1__X2_n, __A09_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9021(net_U9021_Pad1, __A09_1__X2_n, __A09_1__Y2_n, XUY06_n, __A09_1__X2, __A09_1__Y2, GND, __G08_n, CGG, G08, net_U9021_Pad1, XUY06_n, net_U9021_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9022(net_U9022_Pad1, net_U9009_Pad1, net_U9021_Pad1, __A09_1___SUMA2, CO06, __CI07_n, GND, net_U9022_Pad8, __A09_1___SUMA2, __A09_1___SUMB2, RULOG_n, net_U9022_Pad12, G08, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9023(__A09_1___SUMB2, net_U9021_Pad13, net_U9005_Pad12, net_U9023_Pad4, WAG_n, WL06_n, GND, WL08_n, WALSG_n, net_U9023_Pad10, __A09_1___A2_n, CAG, net_U9023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9024(net_U9023_Pad4, net_U9023_Pad10, net_U9022_Pad8, net_U9024_Pad4, CH06, net_U9013_Pad11, GND, net_U9013_Pad13, net_U9024_Pad9, net_U9024_Pad10, net_U9024_Pad11, __A09_1___A2_n, net_U9023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9025(net_U9024_Pad4, RAG_n, __A09_1___A2_n, net_U9024_Pad9, WLG_n, WL06_n, GND, G09_n, G2LSG_n, net_U9024_Pad10, __L06_n, CLG1G, net_U9024_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9026(RLG_n, __L06_n, __A09_1___RL_OUT_2, net_U9026_Pad4, net_U9026_Pad5, net_U9026_Pad6, GND, net_U9026_Pad8, MDT06, R1C, GND, __A09_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9027(net_U9027_Pad1, WQG_n, WL06_n, __A09_1___Q2_n, net_U9027_Pad1, net_U9027_Pad10, GND, __A09_1___Q2_n, CQG, net_U9027_Pad10, RQG_n, __A09_1___Q2_n, net_U9026_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9028(net_U9026_Pad6, RL06_n, net_U9028_Pad3, __A09_1___Z2_n, net_U9026_Pad8, RL06_n, GND, RL06_n, net_U9028_Pad9, G06_n, net_U9018_Pad13, G06_n, net_U9028_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9029(net_U9029_Pad1, WZG_n, WL06_n, net_U9028_Pad3, net_U9029_Pad1, net_U9029_Pad10, GND, __A09_1___Z2_n, CZG, net_U9029_Pad10, RZG_n, __A09_1___Z2_n, net_U9026_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9030(net_U9030_Pad1, WBG_n, WL06_n, __A09_1___B2_n, net_U9030_Pad1, net_U9030_Pad10, GND, __A09_1___B2_n, CBG, net_U9030_Pad10, RBLG_n, __A09_1___B2_n, net_U9030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U9031(net_U9030_Pad13, net_U9031_Pad2, net_U9031_Pad3, net_U9031_Pad4, G06, net_U9028_Pad13, GND, net_U9031_Pad8, GND, XUY10_n, __XUY08_n, net_U9028_Pad9, net_U9031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9032(net_U9031_Pad2, net_U9030_Pad10, RCG_n, net_U9018_Pad11, WL05_n, WG3G_n, GND, WL07_n, WG4G_n, net_U9018_Pad12, L2GDG_n, __L05_n, net_U9031_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9033(net_U9031_Pad4, WG1G_n, WL06_n, G06, G06_n, CGG, GND, RGG_n, G06_n, net_U9031_Pad13, RGG_n, __G08_n, net_U9004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9034(G06_n, GEM06, RL06_n, WL06, WL06, WL06_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9035(net_U9035_Pad1, A2XG_n, __A09_2___A1_n, net_U9035_Pad4, WYLOG_n, WL07_n, GND, WL06_n, WYDG_n, net_U9035_Pad10, __A09_2__Y1_n, CUG, __A09_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9036(MONEX, net_U9035_Pad1, __A09_2__X1_n, CLXC, CUG, __A09_2__X1, GND, __A09_2__Y1_n, net_U9035_Pad4, net_U9035_Pad10, __A09_2__Y1, __A09_2__X1_n, __A09_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9037(net_U9037_Pad1, __A09_2__X1_n, __A09_2__Y1_n, __XUY07_n, __A09_2__X1, __A09_2__Y1, GND, net_U9037_Pad1, __XUY07_n, net_U9037_Pad10, net_U9037_Pad1, __A09_2___SUMA1, __A09_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9038(net_U9038_Pad1, net_U9038_Pad2, __A09_2___SUMA1, __A09_2___SUMB1, RULOG_n, net_U9038_Pad6, GND, net_U9038_Pad8, XUY09_n, __XUY07_n, __CI07_n, net_U9038_Pad12, G07, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9039(__CI07_n, net_U9039_Pad2, G07_n, GEM07, __A09_2___RL1_n, WL07, GND, WL07_n, WL07,  ,  , net_U9039_Pad12, __A09_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9040(__A09_2___SUMB1, net_U9037_Pad10, net_U9039_Pad2, net_U9040_Pad4, WAG_n, WL07_n, GND, WL09_n, WALSG_n, net_U9040_Pad10, __A09_2___A1_n, CAG, net_U9040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9041(net_U9038_Pad8, CO10, net_U9041_Pad3, __A09_2___RL1_n, net_U9041_Pad5, __L07_n, GND, __A09_2___Z1_n, net_U9041_Pad9, __A09_2___RL1_n, net_U9041_Pad11, __A09_2___RL1_n, net_U9041_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1) U9042(net_U9040_Pad4, net_U9040_Pad10, net_U9038_Pad6, net_U9042_Pad4, CH07, net_U9041_Pad3, GND, net_U9041_Pad5, net_U9042_Pad9, net_U9042_Pad10, net_U9042_Pad11, __A09_2___A1_n, net_U9040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9043(net_U9042_Pad4, RAG_n, __A09_2___A1_n, net_U9042_Pad9, WLG_n, WL07_n, GND, G10_n, G2LSG_n, net_U9042_Pad10, __L07_n, CLG1G, net_U9042_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9044(net_U9044_Pad1, __A09_2___SUMA2, __A09_2___SUMA2, __A09_2___SUMB2, RULOG_n, net_U9044_Pad6, GND, __A09_2___RL_OUT_1, RLG_n, __L07_n, GND, CI09_n, __CO08, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9045( ,  ,  , net_U9045_Pad4, WQG_n, WL07_n, GND, net_U9045_Pad4, net_U9045_Pad13, __A09_2___Q1_n, __A09_2___Q1_n, CQG, net_U9045_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9046(net_U9046_Pad1, RQG_n, __A09_2___Q1_n, net_U9046_Pad4, WZG_n, WL07_n, GND, net_U9046_Pad4, net_U9046_Pad13, net_U9041_Pad9, __A09_2___Z1_n, CZG, net_U9046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9047(net_U9047_Pad1, RZG_n, __A09_2___Z1_n, net_U9047_Pad4, WBG_n, WL07_n, GND, net_U9047_Pad4, net_U9047_Pad13, __A09_2___B1_n, __A09_2___B1_n, CBG, net_U9047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9048(net_U9048_Pad1, RBLG_n, __A09_2___B1_n, net_U9048_Pad4, net_U9047_Pad13, RCG_n, GND, WL06_n, WG3G_n, net_U9048_Pad10, WL08_n, WG4G_n, net_U9048_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9049(__A09_2___RL_OUT_1, net_U9046_Pad1, MDT07, R1C, GND, net_U9041_Pad13, GND, net_U9049_Pad8, net_U9048_Pad1, net_U9048_Pad4, net_U9049_Pad11, net_U9041_Pad11, net_U9047_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9050(net_U9031_Pad8, CO10, net_U9049_Pad8, __A09_2___RL1_n, net_U9050_Pad5, G07_n, GND, G07_n, net_U9038_Pad12, __A09_2___RL2_n, net_U9050_Pad11, L08_n, net_U9050_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U9051(net_U9038_Pad1, L2GDG_n, __L06_n, net_U9038_Pad2, WG1G_n, WL07_n, GND, G07_n, CGG, G07, RGG_n, G07_n, net_U9049_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U9052(net_U9050_Pad5, G07ED, SA07, net_U9048_Pad10, net_U9048_Pad13,  , GND,  , GND, SA08, net_U9052_Pad11, net_U9052_Pad12, net_U9052_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9053(net_U9053_Pad1, A2XG_n, __A09_2___A2_n, net_U9053_Pad4, WYLOG_n, WL08_n, GND, WL07_n, WYDG_n, net_U9053_Pad10, __A09_2__Y2_n, CUG, __A09_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9054(MONEX, net_U9053_Pad1, __A09_2__X2_n, CLXC, CUG, __A09_2__X2, GND, __A09_2__Y2_n, net_U9053_Pad4, net_U9053_Pad10, __A09_2__Y2, __A09_2__X2_n, __A09_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9055(net_U9044_Pad1, __A09_2__X2_n, __A09_2__Y2_n, __XUY08_n, __A09_2__X2, __A09_2__Y2, GND,  ,  ,  , net_U9044_Pad1, __XUY08_n, net_U9055_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9056(__A09_2___SUMB2, net_U9055_Pad13, net_U9039_Pad12, net_U9056_Pad4, WAG_n, WL08_n, GND, WL10_n, WALSG_n, net_U9056_Pad10, __A09_2___A2_n, CAG, net_U9056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9057(net_U9056_Pad4, net_U9056_Pad10, net_U9044_Pad6, net_U9057_Pad4, CH08, net_U9050_Pad11, GND, net_U9050_Pad13, net_U9057_Pad9, net_U9057_Pad10, net_U9057_Pad11, __A09_2___A2_n, net_U9056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9058(net_U9057_Pad4, RAG_n, __A09_2___A2_n, net_U9057_Pad9, WLG_n, WL08_n, GND, G11_n, G2LSG_n, net_U9057_Pad10, L08_n, CLG1G, net_U9057_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9059(RLG_n, L08_n, __A09_2___RL_OUT_2, net_U9059_Pad4, net_U9059_Pad5, net_U9059_Pad6, GND, net_U9059_Pad8, MDT08, R1C, GND, __A09_2___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9060(net_U9060_Pad1, WQG_n, WL08_n, __A09_2___Q2_n, net_U9060_Pad1, net_U9060_Pad10, GND, __A09_2___Q2_n, CQG, net_U9060_Pad10, RQG_n, __A09_2___Q2_n, net_U9059_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9061(net_U9059_Pad6, __A09_2___RL2_n, net_U9061_Pad3, __A09_2___Z2_n, net_U9059_Pad8, __A09_2___RL2_n, GND, __A09_2___RL2_n, net_U9004_Pad12, __G08_n, net_U9052_Pad13, __G08_n, net_U9022_Pad12, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9062(net_U9062_Pad1, WZG_n, WL08_n, net_U9061_Pad3, net_U9062_Pad1, net_U9062_Pad10, GND, __A09_2___Z2_n, CZG, net_U9062_Pad10, RZG_n, __A09_2___Z2_n, net_U9059_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9063(net_U9063_Pad1, WBG_n, WL08_n, __A09_2___B2_n, net_U9063_Pad1, net_U9063_Pad10, GND, __A09_2___B2_n, CBG, net_U9063_Pad10, RBLG_n, __A09_2___B2_n, net_U9004_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9064(net_U9004_Pad2, net_U9063_Pad10, RCG_n, net_U9052_Pad11, WL07_n, WG3G_n, GND, WL09_n, WG4G_n, net_U9052_Pad12, L2GDG_n, __L07_n, net_U9022_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9065(__G08_n, GEM08, __A09_2___RL2_n, WL08, WL08, WL08_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U9066(__A09_1___SUMA1, net_U9003_Pad1, XUY05_n, CI05_n, GND,  , GND,  , net_U9021_Pad1, XUY06_n, __A09_1___CI_INTERNAL, GND, __A09_1___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U9067(__A09_2___SUMA1, net_U9037_Pad1, __XUY07_n, __CI07_n, WHOMP,  , GND,  , net_U9044_Pad1, __XUY08_n, __A09_2___CI_INTERNAL, GND, __A09_2___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U9068(RL05_n, MWL05, RL06_n, MWL06, __A09_2___RL1_n, MWL07, GND, MWL08, __A09_2___RL2_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8
endmodule