`timescale 1ns/1ps
`default_nettype none

module four_bit_4(SIM_RST, SIM_CLK, p4VSW, GND, A2XG_n, CAG, CBG, CGG, CLG1G, CLG2G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI13_n, CO14, BXVX, MONEX, XUY01_n, XUY02_n, CH13, CH14, CH16, L12_n, L16_n, G2LSG_n, WL01_n, WL02_n, G01_n, MDT13, MDT14, MDT15, MDT16, SA13, SA14, SA16, RBHG_n, RULOG_n, RUG_n, G16SW_n, WG1G_n, WG2G_n, WG3G_n, WG4G_n, WG5G_n, WYDG_n, WYHIG_n, R1C, US2SG, WL12_n, WHOMPA, Z15_n, Z16_n, A15_n, A16_n, EAC_n, G13, G13_n, G14, G14_n, G15, G15_n, G16, L15_n, RL13_n, RL14_n, RL15_n, RL16_n, SUMA13_n, SUMB13_n, SUMA14_n, SUMB14_n, SUMA15_n, SUMB15_n, SUMA16_n, SUMB16_n, WL13, WL13_n, WL14, WL14_n, WL15, WL15_n, WL16, WL16_n, XUY13_n, XUY14_n, GEM13, GEM14, GEM16, MWL13, MWL14, MWL15, MWL16);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    output wire A15_n;
    output wire A16_n;
    input wire A2XG_n;
    input wire BXVX;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH13;
    input wire CH14;
    input wire CH16;
    input wire CI13_n;
    input wire CLG1G;
    input wire CLG2G;
    input wire CLXC;
    input wire CO14;
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire EAC_n;
    input wire G01_n;
    output wire G13;
    inout wire G13_n; //FPGA#wand
    output wire G14;
    inout wire G14_n; //FPGA#wand
    output wire G15;
    inout wire G15_n; //FPGA#wand
    output wire G16;
    input wire G16SW_n;
    input wire G2LSG_n;
    output wire GEM13;
    output wire GEM14;
    output wire GEM16;
    input wire L12_n;
    inout wire L15_n; //FPGA#wand
    inout wire L16_n; //FPGA#wand
    input wire L2GDG_n;
    input wire MDT13;
    input wire MDT14;
    input wire MDT15;
    input wire MDT16;
    input wire MONEX;
    output wire MWL13; //FPGA#wand
    output wire MWL14; //FPGA#wand
    output wire MWL15; //FPGA#wand
    output wire MWL16; //FPGA#wand
    input wire R1C;
    input wire RAG_n;
    input wire RBHG_n;
    input wire RCG_n;
    input wire RGG_n;
    inout wire RL13_n; //FPGA#wand
    inout wire RL14_n; //FPGA#wand
    inout wire RL15_n; //FPGA#wand
    inout wire RL16_n; //FPGA#wand
    input wire RLG_n;
    input wire RQG_n;
    input wire RUG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA13;
    input wire SA14;
    input wire SA16;
    output wire SUMA13_n;
    output wire SUMA14_n;
    output wire SUMA15_n;
    output wire SUMA16_n;
    output wire SUMB13_n;
    output wire SUMB14_n;
    output wire SUMB15_n;
    output wire SUMB16_n;
    input wire US2SG;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG2G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WG5G_n;
    input wire WHOMPA;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL12_n;
    output wire WL13;
    output wire WL13_n;
    output wire WL14;
    output wire WL14_n;
    output wire WL15;
    output wire WL15_n;
    output wire WL16;
    output wire WL16_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYHIG_n;
    input wire WZG_n;
    input wire XUY01_n;
    input wire XUY02_n;
    output wire XUY13_n;
    output wire XUY14_n;
    inout wire Z15_n; //FPGA#wand
    inout wire Z16_n; //FPGA#wand
    wire __A11_1__X1;
    wire __A11_1__X1_n;
    wire __A11_1__X2;
    wire __A11_1__X2_n;
    wire __A11_1__Y1;
    wire __A11_1__Y1_n;
    wire __A11_1__Y2;
    wire __A11_1__Y2_n;
    wire __A11_1___A1_n;
    wire __A11_1___A2_n;
    wire __A11_1___B1_n;
    wire __A11_1___B2_n;
    wire __A11_1___CI_INTERNAL;
    wire __A11_1___Q1_n;
    wire __A11_1___Q2_n;
    wire __A11_1___RL_OUT_1;
    wire __A11_1___RL_OUT_2;
    wire __A11_1___Z1_n; //FPGA#wand
    wire __A11_1___Z2_n; //FPGA#wand
    wire __A11_2__X1;
    wire __A11_2__X1_n;
    wire __A11_2__X2;
    wire __A11_2__X2_n;
    wire __A11_2__Y1;
    wire __A11_2__Y1_n;
    wire __A11_2__Y2;
    wire __A11_2__Y2_n;
    wire __A11_2___B1_n;
    wire __A11_2___B2_n;
    wire __A11_2___CI_INTERNAL;
    wire __A11_2___CO_OUT; //FPGA#wand
    wire __A11_2___GEM1;
    wire __A11_2___Q1_n;
    wire __A11_2___Q2_n;
    wire __A11_2___RL_OUT_1;
    wire __CI15_n;
    wire __CO16; //FPGA#wand
    wire __G16_n; //FPGA#wand
    wire __L13_n; //FPGA#wand
    wire __L14_n; //FPGA#wand
    wire __RL16;
    wire __XUY15_n;
    wire __XUY16_n;
    wire net_U11001_Pad1;
    wire net_U11001_Pad10;
    wire net_U11001_Pad4;
    wire net_U11003_Pad1;
    wire net_U11003_Pad10;
    wire net_U11004_Pad1;
    wire net_U11004_Pad12;
    wire net_U11004_Pad13;
    wire net_U11004_Pad2;
    wire net_U11004_Pad6;
    wire net_U11004_Pad8;
    wire net_U11005_Pad12;
    wire net_U11005_Pad2;
    wire net_U11006_Pad10;
    wire net_U11006_Pad13;
    wire net_U11006_Pad4;
    wire net_U11007_Pad11;
    wire net_U11007_Pad13;
    wire net_U11007_Pad3;
    wire net_U11007_Pad5;
    wire net_U11007_Pad9;
    wire net_U11008_Pad1;
    wire net_U11008_Pad10;
    wire net_U11008_Pad13;
    wire net_U11008_Pad4;
    wire net_U11009_Pad1;
    wire net_U11009_Pad13;
    wire net_U11009_Pad4;
    wire net_U11010_Pad1;
    wire net_U11010_Pad13;
    wire net_U11010_Pad4;
    wire net_U11011_Pad10;
    wire net_U11011_Pad11;
    wire net_U11011_Pad13;
    wire net_U11011_Pad8;
    wire net_U11011_Pad9;
    wire net_U11012_Pad13;
    wire net_U11012_Pad4;
    wire net_U11013_Pad1;
    wire net_U11013_Pad11;
    wire net_U11013_Pad13;
    wire net_U11013_Pad5;
    wire net_U11013_Pad9;
    wire net_U11014_Pad10;
    wire net_U11014_Pad13;
    wire net_U11016_Pad1;
    wire net_U11016_Pad4;
    wire net_U11018_Pad11;
    wire net_U11018_Pad12;
    wire net_U11018_Pad13;
    wire net_U11019_Pad1;
    wire net_U11019_Pad10;
    wire net_U11019_Pad4;
    wire net_U11021_Pad1;
    wire net_U11021_Pad13;
    wire net_U11022_Pad1;
    wire net_U11022_Pad12;
    wire net_U11022_Pad8;
    wire net_U11023_Pad10;
    wire net_U11023_Pad13;
    wire net_U11023_Pad4;
    wire net_U11024_Pad10;
    wire net_U11024_Pad11;
    wire net_U11024_Pad4;
    wire net_U11024_Pad9;
    wire net_U11026_Pad4;
    wire net_U11026_Pad5;
    wire net_U11026_Pad6;
    wire net_U11026_Pad8;
    wire net_U11027_Pad1;
    wire net_U11027_Pad10;
    wire net_U11028_Pad13;
    wire net_U11028_Pad3;
    wire net_U11028_Pad9;
    wire net_U11029_Pad1;
    wire net_U11029_Pad10;
    wire net_U11030_Pad1;
    wire net_U11030_Pad10;
    wire net_U11030_Pad13;
    wire net_U11031_Pad13;
    wire net_U11031_Pad2;
    wire net_U11031_Pad3;
    wire net_U11031_Pad4;
    wire net_U11031_Pad8;
    wire net_U11035_Pad1;
    wire net_U11035_Pad10;
    wire net_U11035_Pad4;
    wire net_U11037_Pad1;
    wire net_U11037_Pad10;
    wire net_U11038_Pad1;
    wire net_U11038_Pad12;
    wire net_U11038_Pad2;
    wire net_U11038_Pad6;
    wire net_U11038_Pad8;
    wire net_U11039_Pad12;
    wire net_U11039_Pad2;
    wire net_U11040_Pad10;
    wire net_U11040_Pad13;
    wire net_U11040_Pad4;
    wire net_U11041_Pad11;
    wire net_U11041_Pad13;
    wire net_U11041_Pad3;
    wire net_U11041_Pad5;
    wire net_U11041_Pad9;
    wire net_U11042_Pad10;
    wire net_U11042_Pad11;
    wire net_U11042_Pad4;
    wire net_U11042_Pad9;
    wire net_U11044_Pad1;
    wire net_U11044_Pad6;
    wire net_U11045_Pad13;
    wire net_U11045_Pad4;
    wire net_U11046_Pad1;
    wire net_U11046_Pad13;
    wire net_U11046_Pad4;
    wire net_U11047_Pad1;
    wire net_U11047_Pad13;
    wire net_U11047_Pad4;
    wire net_U11048_Pad1;
    wire net_U11048_Pad10;
    wire net_U11048_Pad13;
    wire net_U11048_Pad4;
    wire net_U11049_Pad11;
    wire net_U11049_Pad8;
    wire net_U11050_Pad11;
    wire net_U11050_Pad13;
    wire net_U11050_Pad5;
    wire net_U11052_Pad11;
    wire net_U11052_Pad12;
    wire net_U11052_Pad13;
    wire net_U11053_Pad1;
    wire net_U11053_Pad10;
    wire net_U11053_Pad4;
    wire net_U11055_Pad13;
    wire net_U11056_Pad10;
    wire net_U11056_Pad13;
    wire net_U11056_Pad4;
    wire net_U11057_Pad10;
    wire net_U11057_Pad11;
    wire net_U11057_Pad4;
    wire net_U11057_Pad9;
    wire net_U11059_Pad4;
    wire net_U11059_Pad5;
    wire net_U11059_Pad6;
    wire net_U11059_Pad8;
    wire net_U11060_Pad1;
    wire net_U11060_Pad10;
    wire net_U11061_Pad3;
    wire net_U11062_Pad1;
    wire net_U11062_Pad10;
    wire net_U11063_Pad1;
    wire net_U11063_Pad10;

    pullup R11001(__CO16);
    pullup R11002(RL13_n);
    pullup R11003(__L13_n);
    pullup R11005(__A11_1___Z1_n);
    pullup R11006(G13_n);
    pullup R11007(RL14_n);
    pullup R11008(__L14_n);
    pullup R11009(__A11_1___Z2_n);
    pullup R11010(G14_n);
    pullup R11011(__A11_2___CO_OUT);
    pullup R11012(RL15_n);
    pullup R11013(L15_n);
    pullup R11015(Z15_n);
    pullup R11016(G15_n);
    pullup R11017(RL16_n);
    pullup R11018(L16_n);
    pullup R11019(Z16_n);
    pullup R11020(__G16_n);
    U74HC02 U11001(net_U11001_Pad1, A2XG_n, __A11_1___A1_n, net_U11001_Pad4, WYHIG_n, WL13_n, GND, WL12_n, WYDG_n, net_U11001_Pad10, __A11_1__Y1_n, CUG, __A11_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11002(MONEX, net_U11001_Pad1, __A11_1__X1_n, CLXC, CUG, __A11_1__X1, GND, __A11_1__Y1_n, net_U11001_Pad4, net_U11001_Pad10, __A11_1__Y1, __A11_1__X1_n, __A11_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11003(net_U11003_Pad1, __A11_1__X1_n, __A11_1__Y1_n, XUY13_n, __A11_1__X1, __A11_1__Y1, GND, net_U11003_Pad1, XUY13_n, net_U11003_Pad10, net_U11003_Pad1, SUMA13_n, __A11_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11004(net_U11004_Pad1, net_U11004_Pad2, SUMA13_n, SUMB13_n, RULOG_n, net_U11004_Pad6, GND, net_U11004_Pad8, __XUY15_n, XUY13_n, CI13_n, net_U11004_Pad12, net_U11004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11005(CI13_n, net_U11005_Pad2, G13_n, GEM13, RL13_n, WL13, GND, WL13_n, WL13,  ,  , net_U11005_Pad12, __A11_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11006(SUMB13_n, net_U11003_Pad10, net_U11005_Pad2, net_U11006_Pad4, WAG_n, WL13_n, GND, WL15_n, WALSG_n, net_U11006_Pad10, __A11_1___A1_n, CAG, net_U11006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11007(net_U11004_Pad8, __CO16, net_U11007_Pad3, RL13_n, net_U11007_Pad5, __L13_n, GND, __A11_1___Z1_n, net_U11007_Pad9, RL13_n, net_U11007_Pad11, RL13_n, net_U11007_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U11008(net_U11008_Pad1, RAG_n, __A11_1___A1_n, net_U11008_Pad4, WLG_n, WL13_n, GND, WL01_n, WALSG_n, net_U11008_Pad10, __L13_n, CLG2G, net_U11008_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11009(net_U11009_Pad1, WG2G_n, WL16_n, net_U11009_Pad4, WQG_n, WL13_n, GND, net_U11009_Pad4, net_U11009_Pad13, __A11_1___Q1_n, __A11_1___Q1_n, CQG, net_U11009_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11010(net_U11010_Pad1, RQG_n, __A11_1___Q1_n, net_U11010_Pad4, WZG_n, WL13_n, GND, net_U11010_Pad4, net_U11010_Pad13, net_U11007_Pad9, __A11_1___Z1_n, CZG, net_U11010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11011(__A11_1___RL_OUT_1, net_U11010_Pad1, MDT13, R1C, GND, net_U11007_Pad13, GND, net_U11011_Pad8, net_U11011_Pad9, net_U11011_Pad10, net_U11011_Pad11, net_U11007_Pad11, net_U11011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11012(net_U11011_Pad13, RZG_n, __A11_1___Z1_n, net_U11012_Pad4, WBG_n, WL13_n, GND, net_U11012_Pad4, net_U11012_Pad13, __A11_1___B1_n, __A11_1___B1_n, CBG, net_U11012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11013(net_U11013_Pad1, __CO16, net_U11011_Pad8, RL13_n, net_U11013_Pad5, G13_n, GND, G13_n, net_U11013_Pad9, RL14_n, net_U11013_Pad11, __L14_n, net_U11013_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U11014(net_U11011_Pad9, RBHG_n, __A11_1___B1_n, net_U11011_Pad10, net_U11012_Pad13, RCG_n, GND, WL12_n, WG3G_n, net_U11014_Pad10, WL14_n, WG4G_n, net_U11014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11015(net_U11006_Pad4, net_U11006_Pad10, net_U11004_Pad6, net_U11008_Pad1, CH13, net_U11007_Pad3, GND, net_U11007_Pad5, net_U11008_Pad4, net_U11008_Pad10, net_U11008_Pad13, __A11_1___A1_n, net_U11006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11016(net_U11016_Pad1, L2GDG_n, L12_n, net_U11016_Pad4, WG1G_n, WL13_n, GND, G13_n, CGG, G13, RGG_n, G13_n, net_U11011_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11017(net_U11016_Pad1, net_U11016_Pad4, GND, __XUY16_n, XUY14_n, net_U11013_Pad1, GND, __A11_1___RL_OUT_1, RLG_n, __L13_n, GND, net_U11013_Pad9, G13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U11018(net_U11013_Pad5, GND, SA13, net_U11014_Pad10, net_U11014_Pad13,  , GND,  , GND, SA14, net_U11018_Pad11, net_U11018_Pad12, net_U11018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11019(net_U11019_Pad1, A2XG_n, __A11_1___A2_n, net_U11019_Pad4, WYHIG_n, WL14_n, GND, WL13_n, WYDG_n, net_U11019_Pad10, __A11_1__Y2_n, CUG, __A11_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11020(MONEX, net_U11019_Pad1, __A11_1__X2_n, CLXC, CUG, __A11_1__X2, GND, __A11_1__Y2_n, net_U11019_Pad4, net_U11019_Pad10, __A11_1__Y2, __A11_1__X2_n, __A11_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11021(net_U11021_Pad1, __A11_1__X2_n, __A11_1__Y2_n, XUY14_n, __A11_1__X2, __A11_1__Y2, GND, __G16_n, CGG, G16, net_U11021_Pad1, XUY14_n, net_U11021_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11022(net_U11022_Pad1, net_U11009_Pad1, net_U11021_Pad1, SUMA14_n, CO14, __CI15_n, GND, net_U11022_Pad8, SUMA14_n, SUMB14_n, RULOG_n, net_U11022_Pad12, G16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11023(SUMB14_n, net_U11021_Pad13, net_U11005_Pad12, net_U11023_Pad4, WAG_n, WL14_n, GND, WL16_n, WALSG_n, net_U11023_Pad10, __A11_1___A2_n, CAG, net_U11023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11024(net_U11023_Pad4, net_U11023_Pad10, net_U11022_Pad8, net_U11024_Pad4, CH14, net_U11013_Pad11, GND, net_U11013_Pad13, net_U11024_Pad9, net_U11024_Pad10, net_U11024_Pad11, __A11_1___A2_n, net_U11023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11025(net_U11024_Pad4, RAG_n, __A11_1___A2_n, net_U11024_Pad9, WLG_n, WL14_n, GND, WL02_n, WALSG_n, net_U11024_Pad10, __L14_n, CLG2G, net_U11024_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11026(RLG_n, __L14_n, __A11_1___RL_OUT_2, net_U11026_Pad4, net_U11026_Pad5, net_U11026_Pad6, GND, net_U11026_Pad8, MDT14, R1C, GND, __A11_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11027(net_U11027_Pad1, WQG_n, WL14_n, __A11_1___Q2_n, net_U11027_Pad1, net_U11027_Pad10, GND, __A11_1___Q2_n, CQG, net_U11027_Pad10, RQG_n, __A11_1___Q2_n, net_U11026_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11028(net_U11026_Pad6, RL14_n, net_U11028_Pad3, __A11_1___Z2_n, net_U11026_Pad8, RL14_n, GND, RL14_n, net_U11028_Pad9, G14_n, net_U11018_Pad13, G14_n, net_U11028_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11029(net_U11029_Pad1, WZG_n, WL14_n, net_U11028_Pad3, net_U11029_Pad1, net_U11029_Pad10, GND, __A11_1___Z2_n, CZG, net_U11029_Pad10, RZG_n, __A11_1___Z2_n, net_U11026_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11030(net_U11030_Pad1, WBG_n, WL14_n, __A11_1___B2_n, net_U11030_Pad1, net_U11030_Pad10, GND, __A11_1___B2_n, CBG, net_U11030_Pad10, RBHG_n, __A11_1___B2_n, net_U11030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U11031(net_U11030_Pad13, net_U11031_Pad2, net_U11031_Pad3, net_U11031_Pad4, G14, net_U11028_Pad13, GND, net_U11031_Pad8, GND, XUY02_n, __XUY16_n, net_U11028_Pad9, net_U11031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11032(net_U11031_Pad2, net_U11030_Pad10, RCG_n, net_U11018_Pad11, WL13_n, WG3G_n, GND, WL16_n, WG4G_n, net_U11018_Pad12, L2GDG_n, __L13_n, net_U11031_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11033(net_U11031_Pad4, WG1G_n, WL14_n, G14, G14_n, CGG, GND, RGG_n, G14_n, net_U11031_Pad13, RGG_n, __G16_n, net_U11004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11034(G14_n, GEM14, RL14_n, WL14, WL14, WL14_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11035(net_U11035_Pad1, A2XG_n, A15_n, net_U11035_Pad4, WYHIG_n, WL15_n, GND, WL14_n, WYDG_n, net_U11035_Pad10, __A11_2__Y1_n, CUG, __A11_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11036(BXVX, net_U11035_Pad1, __A11_2__X1_n, CLXC, CUG, __A11_2__X1, GND, __A11_2__Y1_n, net_U11035_Pad4, net_U11035_Pad10, __A11_2__Y1, __A11_2__X1_n, __A11_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11037(net_U11037_Pad1, __A11_2__X1_n, __A11_2__Y1_n, __XUY15_n, __A11_2__X1, __A11_2__Y1, GND, net_U11037_Pad1, __XUY15_n, net_U11037_Pad10, net_U11037_Pad1, SUMA15_n, __A11_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11038(net_U11038_Pad1, net_U11038_Pad2, SUMA15_n, SUMB15_n, RULOG_n, net_U11038_Pad6, GND, net_U11038_Pad8, XUY01_n, __XUY15_n, __CI15_n, net_U11038_Pad12, G15, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11039(__CI15_n, net_U11039_Pad2, G15_n, __A11_2___GEM1, RL15_n, WL15, GND, WL15_n, WL15,  ,  , net_U11039_Pad12, __A11_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11040(SUMB15_n, net_U11037_Pad10, net_U11039_Pad2, net_U11040_Pad4, WAG_n, WL15_n, GND, G16SW_n, WALSG_n, net_U11040_Pad10, A15_n, CAG, net_U11040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11041(net_U11038_Pad8, __A11_2___CO_OUT, net_U11041_Pad3, RL15_n, net_U11041_Pad5, L15_n, GND, Z15_n, net_U11041_Pad9, RL15_n, net_U11041_Pad11, RL15_n, net_U11041_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1) U11042(net_U11040_Pad4, net_U11040_Pad10, net_U11038_Pad6, net_U11042_Pad4, CH16, net_U11041_Pad3, GND, net_U11041_Pad5, net_U11042_Pad9, net_U11042_Pad10, net_U11042_Pad11, A15_n, net_U11040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11043(net_U11042_Pad4, RAG_n, A15_n, net_U11042_Pad9, WLG_n, WL15_n, GND, G01_n, G2LSG_n, net_U11042_Pad10, L15_n, CLG1G, net_U11042_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11044(net_U11044_Pad1, SUMA16_n, SUMA16_n, SUMB16_n, RUG_n, net_U11044_Pad6, GND, __A11_2___RL_OUT_1, RLG_n, L15_n, p4VSW, EAC_n, __CO16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11045( ,  ,  , net_U11045_Pad4, WQG_n, WL15_n, GND, net_U11045_Pad4, net_U11045_Pad13, __A11_2___Q1_n, __A11_2___Q1_n, CQG, net_U11045_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11046(net_U11046_Pad1, RQG_n, __A11_2___Q1_n, net_U11046_Pad4, WZG_n, WL15_n, GND, net_U11046_Pad4, net_U11046_Pad13, net_U11041_Pad9, Z15_n, CZG, net_U11046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11047(net_U11047_Pad1, RZG_n, Z15_n, net_U11047_Pad4, WBG_n, WL15_n, GND, net_U11047_Pad4, net_U11047_Pad13, __A11_2___B1_n, __A11_2___B1_n, CBG, net_U11047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11048(net_U11048_Pad1, RBHG_n, __A11_2___B1_n, net_U11048_Pad4, net_U11047_Pad13, RCG_n, GND, GND, p4VSW, net_U11048_Pad10, GND, p4VSW, net_U11048_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11049(__A11_2___RL_OUT_1, net_U11046_Pad1, MDT15, R1C, __RL16, net_U11041_Pad13, GND, net_U11049_Pad8, net_U11048_Pad1, net_U11048_Pad4, net_U11049_Pad11, net_U11041_Pad11, net_U11047_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11050(net_U11031_Pad8, __A11_2___CO_OUT, net_U11049_Pad8, RL15_n, net_U11050_Pad5, G15_n, GND, G15_n, net_U11038_Pad12, RL16_n, net_U11050_Pad11, L16_n, net_U11050_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U11051(net_U11038_Pad1, L2GDG_n, __L14_n, net_U11038_Pad2, WG1G_n, WL15_n, GND, G15_n, CGG, G15, RGG_n, G15_n, net_U11049_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U11052(net_U11050_Pad5, GND, SA16, net_U11048_Pad10, net_U11048_Pad13,  , GND,  , GND, SA16, net_U11052_Pad11, net_U11052_Pad12, net_U11052_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11053(net_U11053_Pad1, A2XG_n, A16_n, net_U11053_Pad4, WYHIG_n, WL16_n, GND, WL16_n, WYDG_n, net_U11053_Pad10, __A11_2__Y2_n, CUG, __A11_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11054(MONEX, net_U11053_Pad1, __A11_2__X2_n, CLXC, CUG, __A11_2__X2, GND, __A11_2__Y2_n, net_U11053_Pad4, net_U11053_Pad10, __A11_2__Y2, __A11_2__X2_n, __A11_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11055(net_U11044_Pad1, __A11_2__X2_n, __A11_2__Y2_n, __XUY16_n, __A11_2__X2, __A11_2__Y2, GND,  ,  ,  , net_U11044_Pad1, __XUY16_n, net_U11055_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11056(SUMB16_n, net_U11055_Pad13, net_U11039_Pad12, net_U11056_Pad4, WAG_n, WL16_n, GND, G16SW_n, WALSG_n, net_U11056_Pad10, A16_n, CAG, net_U11056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11057(net_U11056_Pad4, net_U11056_Pad10, net_U11044_Pad6, net_U11057_Pad4, CH16, net_U11050_Pad11, GND, net_U11050_Pad13, net_U11057_Pad9, net_U11057_Pad10, net_U11057_Pad11, A16_n, net_U11056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11058(net_U11057_Pad4, RAG_n, A16_n, net_U11057_Pad9, WLG_n, WL16_n, GND, __G16_n, G2LSG_n, net_U11057_Pad10, L16_n, CLG1G, net_U11057_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11059(RLG_n, L16_n, __RL16, net_U11059_Pad4, net_U11059_Pad5, net_U11059_Pad6, GND, net_U11059_Pad8, MDT16, R1C, US2SG, __RL16, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11060(net_U11060_Pad1, WQG_n, WL16_n, __A11_2___Q2_n, net_U11060_Pad1, net_U11060_Pad10, GND, __A11_2___Q2_n, CQG, net_U11060_Pad10, RQG_n, __A11_2___Q2_n, net_U11059_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11061(net_U11059_Pad6, RL16_n, net_U11061_Pad3, Z16_n, net_U11059_Pad8, RL16_n, GND, RL16_n, net_U11004_Pad12, __G16_n, net_U11052_Pad13, __G16_n, net_U11022_Pad12, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11062(net_U11062_Pad1, WZG_n, WL16_n, net_U11061_Pad3, net_U11062_Pad1, net_U11062_Pad10, GND, Z16_n, CZG, net_U11062_Pad10, RZG_n, Z16_n, net_U11059_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11063(net_U11063_Pad1, WBG_n, WL16_n, __A11_2___B2_n, net_U11063_Pad1, net_U11063_Pad10, GND, __A11_2___B2_n, CBG, net_U11063_Pad10, RBHG_n, __A11_2___B2_n, net_U11004_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11064(net_U11004_Pad2, net_U11063_Pad10, RCG_n, net_U11052_Pad11, WL14_n, WG3G_n, GND, WL01_n, WG5G_n, net_U11052_Pad12, L2GDG_n, L16_n, net_U11022_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11065(__G16_n, GEM16, RL16_n, WL16, WL16, WL16_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U11066(SUMA13_n, net_U11003_Pad1, XUY13_n, CI13_n, GND,  , GND,  , net_U11021_Pad1, XUY14_n, __A11_1___CI_INTERNAL, GND, SUMA14_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U11067(SUMA15_n, net_U11037_Pad1, __XUY15_n, __CI15_n, GND,  , GND,  , net_U11044_Pad1, __XUY16_n, __A11_2___CI_INTERNAL, WHOMPA, SUMA16_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U11068(RL13_n, MWL13, RL14_n, MWL14, RL15_n, MWL15, GND, MWL16, RL16_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8
endmodule