`timescale 1ns/1ps
`default_nettype none

module scaler(SIM_RST, SIM_CLK, p4VDC, GND, FS01_n, RCHAT_n, RCHBT_n, FS02, F02B, FS03, F03B, FS04, F04A, F04B, FS05, FS05_n, F05A_n, F05B_n, FS06, F06B, FS07A, FS07_n, F07A, F07B, F07B_n, FS08, F08B, FS09, FS09_n, F09A, F09B, F09B_n, FS10, F10A, F10A_n, F10B, F12B, FS13, FS14, F14B, FS16, FS17, F17A, F17B, F18A, F18B, CHAT01, CHAT02, CHAT03, CHAT04, CHAT05, CHAT06, CHAT07, CHAT08, CHAT09, CHAT10, CHAT11, CHAT12, CHAT13, CHAT14, CHBT01, CHBT02, CHBT03, CHBT04, CHBT05, CHBT06, CHBT07, CHBT08, CHBT09, CHBT10, CHBT11, CHBT12, CHBT13, CHBT14);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VDC;
    input wire GND;
    output wire CHAT01;
    output wire CHAT02;
    output wire CHAT03;
    output wire CHAT04;
    output wire CHAT05;
    output wire CHAT06;
    output wire CHAT07;
    output wire CHAT08;
    output wire CHAT09;
    output wire CHAT10;
    output wire CHAT11;
    output wire CHAT12;
    output wire CHAT13;
    output wire CHAT14;
    output wire CHBT01;
    output wire CHBT02;
    output wire CHBT03;
    output wire CHBT04;
    output wire CHBT05;
    output wire CHBT06;
    output wire CHBT07;
    output wire CHBT08;
    output wire CHBT09;
    output wire CHBT10;
    output wire CHBT11;
    output wire CHBT12;
    output wire CHBT13;
    output wire CHBT14;
    output wire F02B;
    output wire F03B;
    output wire F04A;
    output wire F04B;
    output wire F05A_n;
    output wire F05B_n;
    output wire F06B;
    output wire F07A;
    output wire F07B;
    output wire F07B_n;
    output wire F08B;
    output wire F09A;
    output wire F09B;
    output wire F09B_n;
    output wire F10A;
    output wire F10A_n;
    output wire F10B;
    output wire F12B;
    output wire F14B;
    output wire F17A;
    output wire F17B;
    output wire F18A;
    output wire F18B;
    input wire FS01_n;
    output wire FS02;
    output wire FS03;
    output wire FS04;
    output wire FS05;
    output wire FS05_n;
    output wire FS06;
    output wire FS07A;
    output wire FS07_n;
    output wire FS08;
    output wire FS09;
    output wire FS09_n;
    output wire FS10;
    output wire FS13;
    output wire FS14;
    output wire FS16;
    output wire FS17;
    input wire RCHAT_n;
    input wire RCHBT_n;
    wire __A01_1__F02A;
    wire __A01_1__F03A;
    wire __A01_1__F05A;
    wire __A01_1__F05B;
    wire __A01_1__F06A;
    wire __A01_1__F08A;
    wire __A01_1__F11A;
    wire __A01_1__F11B;
    wire __A01_1__F12A;
    wire __A01_1__F13A;
    wire __A01_1__F13B;
    wire __A01_1__F14A;
    wire __A01_1__F15A;
    wire __A01_1__F15B;
    wire __A01_1__F16A;
    wire __A01_1__F16B;
    wire __A01_1__FS02A;
    wire __A01_1__FS03A;
    wire __A01_1__FS04A;
    wire __A01_1__FS05A;
    wire __A01_1__FS07;
    wire __A01_1__FS11;
    wire __A01_1__FS12;
    wire __A01_1__FS15;
    wire __A01_1__scaler_s10__FS_n;
    wire __A01_1__scaler_s11__FS_n;
    wire __A01_1__scaler_s12__FS_n;
    wire __A01_1__scaler_s13__FS_n;
    wire __A01_1__scaler_s14__FS_n;
    wire __A01_1__scaler_s15__FS_n;
    wire __A01_1__scaler_s16__FS_n;
    wire __A01_1__scaler_s17__FS_n;
    wire __A01_1__scaler_s2__FS_n;
    wire __A01_1__scaler_s3__FS_n;
    wire __A01_1__scaler_s4__FS_n;
    wire __A01_1__scaler_s5__FS_n;
    wire __A01_1__scaler_s6__FS_n;
    wire __A01_1__scaler_s7__FS_n;
    wire __A01_1__scaler_s8__FS_n;
    wire __A01_1__scaler_s9__FS_n;
    wire __A01_2__F19A;
    wire __A01_2__F19B;
    wire __A01_2__F20A;
    wire __A01_2__F20B;
    wire __A01_2__F21A;
    wire __A01_2__F21B;
    wire __A01_2__F22A;
    wire __A01_2__F22B;
    wire __A01_2__F23A;
    wire __A01_2__F23B;
    wire __A01_2__F24A;
    wire __A01_2__F24B;
    wire __A01_2__F25A;
    wire __A01_2__F25B;
    wire __A01_2__F26A;
    wire __A01_2__F26B;
    wire __A01_2__F27A;
    wire __A01_2__F27B;
    wire __A01_2__F28A;
    wire __A01_2__F28B;
    wire __A01_2__F29A;
    wire __A01_2__F29B;
    wire __A01_2__F30A;
    wire __A01_2__F30B;
    wire __A01_2__F31A;
    wire __A01_2__F31B;
    wire __A01_2__F32A;
    wire __A01_2__F32B;
    wire __A01_2__F33A;
    wire __A01_2__F33B;
    wire __A01_2__FS18;
    wire __A01_2__FS19;
    wire __A01_2__FS20;
    wire __A01_2__FS21;
    wire __A01_2__FS22;
    wire __A01_2__FS23;
    wire __A01_2__FS24;
    wire __A01_2__FS25;
    wire __A01_2__FS26;
    wire __A01_2__FS27;
    wire __A01_2__FS28;
    wire __A01_2__FS29;
    wire __A01_2__FS30;
    wire __A01_2__FS31;
    wire __A01_2__FS32;
    wire __A01_2__FS33;
    wire __A01_2__scaler_s18__FS_n;
    wire __A01_2__scaler_s19__FS_n;
    wire __A01_2__scaler_s20__FS_n;
    wire __A01_2__scaler_s21__FS_n;
    wire __A01_2__scaler_s22__FS_n;
    wire __A01_2__scaler_s23__FS_n;
    wire __A01_2__scaler_s24__FS_n;
    wire __A01_2__scaler_s25__FS_n;
    wire __A01_2__scaler_s26__FS_n;
    wire __A01_2__scaler_s27__FS_n;
    wire __A01_2__scaler_s28__FS_n;
    wire __A01_2__scaler_s29__FS_n;
    wire __A01_2__scaler_s30__FS_n;
    wire __A01_2__scaler_s31__FS_n;
    wire __A01_2__scaler_s32__FS_n;
    wire __A01_2__scaler_s33__FS_n;
    wire net_U1101_Pad12;
    wire net_U1101_Pad3;
    wire net_U1102_Pad11;
    wire net_U1102_Pad8;
    wire net_U1104_Pad5;
    wire net_U1104_Pad6;
    wire net_U1106_Pad12;
    wire net_U1106_Pad3;
    wire net_U1107_Pad11;
    wire net_U1107_Pad8;
    wire net_U1109_Pad5;
    wire net_U1109_Pad6;
    wire net_U1111_Pad12;
    wire net_U1111_Pad3;
    wire net_U1112_Pad11;
    wire net_U1112_Pad8;
    wire net_U1114_Pad5;
    wire net_U1114_Pad6;
    wire net_U1116_Pad12;
    wire net_U1116_Pad3;
    wire net_U1117_Pad11;
    wire net_U1117_Pad8;
    wire net_U1119_Pad5;
    wire net_U1119_Pad6;
    wire net_U1121_Pad12;
    wire net_U1121_Pad3;
    wire net_U1122_Pad11;
    wire net_U1122_Pad8;
    wire net_U1124_Pad5;
    wire net_U1124_Pad6;
    wire net_U1126_Pad12;
    wire net_U1126_Pad3;
    wire net_U1132_Pad12;
    wire net_U1132_Pad3;
    wire net_U1133_Pad11;
    wire net_U1133_Pad8;
    wire net_U1135_Pad5;
    wire net_U1135_Pad6;
    wire net_U1137_Pad12;
    wire net_U1137_Pad3;
    wire net_U1138_Pad11;
    wire net_U1138_Pad8;
    wire net_U1140_Pad5;
    wire net_U1140_Pad6;
    wire net_U1142_Pad12;
    wire net_U1142_Pad3;
    wire net_U1143_Pad11;
    wire net_U1143_Pad8;
    wire net_U1145_Pad5;
    wire net_U1145_Pad6;
    wire net_U1147_Pad12;
    wire net_U1147_Pad3;
    wire net_U1148_Pad11;
    wire net_U1148_Pad8;
    wire net_U1150_Pad5;
    wire net_U1150_Pad6;
    wire net_U1152_Pad12;
    wire net_U1152_Pad3;
    wire net_U1153_Pad11;
    wire net_U1153_Pad8;
    wire net_U1155_Pad5;
    wire net_U1155_Pad6;
    wire net_U1157_Pad12;
    wire net_U1157_Pad3;

    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1101(__A01_1__F02A, __A01_1__scaler_s2__FS_n, net_U1101_Pad3, F02B, net_U1101_Pad12, FS02, GND, net_U1101_Pad3, FS02, __A01_1__scaler_s2__FS_n, __A01_1__scaler_s2__FS_n, net_U1101_Pad12, FS02, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1102(__A01_1__F02A, FS01_n, net_U1101_Pad3, FS01_n, F02B, net_U1101_Pad12, GND, net_U1102_Pad8, __A01_1__F03A, __A01_1__F02A, net_U1102_Pad11, net_U1101_Pad3, net_U1101_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1103(__A01_1__F03A, __A01_1__scaler_s3__FS_n, net_U1102_Pad8, F03B, net_U1102_Pad11, FS03, GND, net_U1102_Pad8, FS03, __A01_1__scaler_s3__FS_n, __A01_1__scaler_s3__FS_n, net_U1102_Pad11, FS03, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1104(net_U1102_Pad8, __A01_1__F02A, F04A, __A01_1__F03A, net_U1104_Pad5, net_U1104_Pad6, GND, net_U1104_Pad5, net_U1104_Pad6, __A01_1__F03A, F04B, net_U1102_Pad11, F03B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1105(F04A, __A01_1__scaler_s4__FS_n, net_U1104_Pad6, F04B, net_U1104_Pad5, FS04, GND, net_U1104_Pad6, FS04, __A01_1__scaler_s4__FS_n, __A01_1__scaler_s4__FS_n, net_U1104_Pad5, FS04, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1106(__A01_1__F05A, __A01_1__scaler_s5__FS_n, net_U1106_Pad3, __A01_1__F05B, net_U1106_Pad12, FS05, GND, net_U1106_Pad3, FS05, __A01_1__scaler_s5__FS_n, __A01_1__scaler_s5__FS_n, net_U1106_Pad12, FS05, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1107(__A01_1__F05A, F04A, net_U1106_Pad3, F04A, __A01_1__F05B, net_U1106_Pad12, GND, net_U1107_Pad8, __A01_1__F06A, __A01_1__F05A, net_U1107_Pad11, net_U1106_Pad3, net_U1106_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1108(__A01_1__F06A, __A01_1__scaler_s6__FS_n, net_U1107_Pad8, F06B, net_U1107_Pad11, FS06, GND, net_U1107_Pad8, FS06, __A01_1__scaler_s6__FS_n, __A01_1__scaler_s6__FS_n, net_U1107_Pad11, FS06, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1109(net_U1107_Pad8, __A01_1__F05A, F07A, __A01_1__F06A, net_U1109_Pad5, net_U1109_Pad6, GND, net_U1109_Pad5, net_U1109_Pad6, __A01_1__F06A, F07B, net_U1107_Pad11, F06B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1110(F07A, __A01_1__scaler_s7__FS_n, net_U1109_Pad6, F07B, net_U1109_Pad5, __A01_1__FS07, GND, net_U1109_Pad6, __A01_1__FS07, __A01_1__scaler_s7__FS_n, __A01_1__scaler_s7__FS_n, net_U1109_Pad5, __A01_1__FS07, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1111(__A01_1__F08A, __A01_1__scaler_s8__FS_n, net_U1111_Pad3, F08B, net_U1111_Pad12, FS08, GND, net_U1111_Pad3, FS08, __A01_1__scaler_s8__FS_n, __A01_1__scaler_s8__FS_n, net_U1111_Pad12, FS08, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1112(__A01_1__F08A, F07A, net_U1111_Pad3, F07A, F08B, net_U1111_Pad12, GND, net_U1112_Pad8, F09A, __A01_1__F08A, net_U1112_Pad11, net_U1111_Pad3, net_U1111_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1113(F09A, __A01_1__scaler_s9__FS_n, net_U1112_Pad8, F09B, net_U1112_Pad11, FS09, GND, net_U1112_Pad8, FS09, __A01_1__scaler_s9__FS_n, __A01_1__scaler_s9__FS_n, net_U1112_Pad11, FS09, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1114(net_U1112_Pad8, __A01_1__F08A, F10A, F09A, net_U1114_Pad5, net_U1114_Pad6, GND, net_U1114_Pad5, net_U1114_Pad6, F09A, F10B, net_U1112_Pad11, F09B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1115(F10A, __A01_1__scaler_s10__FS_n, net_U1114_Pad6, F10B, net_U1114_Pad5, FS10, GND, net_U1114_Pad6, FS10, __A01_1__scaler_s10__FS_n, __A01_1__scaler_s10__FS_n, net_U1114_Pad5, FS10, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1116(__A01_1__F11A, __A01_1__scaler_s11__FS_n, net_U1116_Pad3, __A01_1__F11B, net_U1116_Pad12, __A01_1__FS11, GND, net_U1116_Pad3, __A01_1__FS11, __A01_1__scaler_s11__FS_n, __A01_1__scaler_s11__FS_n, net_U1116_Pad12, __A01_1__FS11, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1117(__A01_1__F11A, F10A, net_U1116_Pad3, F10A, __A01_1__F11B, net_U1116_Pad12, GND, net_U1117_Pad8, __A01_1__F12A, __A01_1__F11A, net_U1117_Pad11, net_U1116_Pad3, net_U1116_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1118(__A01_1__F12A, __A01_1__scaler_s12__FS_n, net_U1117_Pad8, F12B, net_U1117_Pad11, __A01_1__FS12, GND, net_U1117_Pad8, __A01_1__FS12, __A01_1__scaler_s12__FS_n, __A01_1__scaler_s12__FS_n, net_U1117_Pad11, __A01_1__FS12, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1119(net_U1117_Pad8, __A01_1__F11A, __A01_1__F13A, __A01_1__F12A, net_U1119_Pad5, net_U1119_Pad6, GND, net_U1119_Pad5, net_U1119_Pad6, __A01_1__F12A, __A01_1__F13B, net_U1117_Pad11, F12B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1120(__A01_1__F13A, __A01_1__scaler_s13__FS_n, net_U1119_Pad6, __A01_1__F13B, net_U1119_Pad5, FS13, GND, net_U1119_Pad6, FS13, __A01_1__scaler_s13__FS_n, __A01_1__scaler_s13__FS_n, net_U1119_Pad5, FS13, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1121(__A01_1__F14A, __A01_1__scaler_s14__FS_n, net_U1121_Pad3, F14B, net_U1121_Pad12, FS14, GND, net_U1121_Pad3, FS14, __A01_1__scaler_s14__FS_n, __A01_1__scaler_s14__FS_n, net_U1121_Pad12, FS14, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1122(__A01_1__F14A, __A01_1__F13A, net_U1121_Pad3, __A01_1__F13A, F14B, net_U1121_Pad12, GND, net_U1122_Pad8, __A01_1__F15A, __A01_1__F14A, net_U1122_Pad11, net_U1121_Pad3, net_U1121_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1123(__A01_1__F15A, __A01_1__scaler_s15__FS_n, net_U1122_Pad8, __A01_1__F15B, net_U1122_Pad11, __A01_1__FS15, GND, net_U1122_Pad8, __A01_1__FS15, __A01_1__scaler_s15__FS_n, __A01_1__scaler_s15__FS_n, net_U1122_Pad11, __A01_1__FS15, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1124(net_U1122_Pad8, __A01_1__F14A, __A01_1__F16A, __A01_1__F15A, net_U1124_Pad5, net_U1124_Pad6, GND, net_U1124_Pad5, net_U1124_Pad6, __A01_1__F15A, __A01_1__F16B, net_U1122_Pad11, __A01_1__F15B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1125(__A01_1__F16A, __A01_1__scaler_s16__FS_n, net_U1124_Pad6, __A01_1__F16B, net_U1124_Pad5, FS16, GND, net_U1124_Pad6, FS16, __A01_1__scaler_s16__FS_n, __A01_1__scaler_s16__FS_n, net_U1124_Pad5, FS16, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1126(F17A, __A01_1__scaler_s17__FS_n, net_U1126_Pad3, F17B, net_U1126_Pad12, FS17, GND, net_U1126_Pad3, FS17, __A01_1__scaler_s17__FS_n, __A01_1__scaler_s17__FS_n, net_U1126_Pad12, FS17, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1127(F17A, __A01_1__F16A, net_U1126_Pad3, __A01_1__F16A, F17B, net_U1126_Pad12, GND,  ,  ,  ,  , net_U1126_Pad3, net_U1126_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U1128(__A01_1__scaler_s2__FS_n, __A01_1__FS02A, __A01_1__scaler_s3__FS_n, __A01_1__FS03A, __A01_1__scaler_s4__FS_n, __A01_1__FS04A, GND, __A01_1__FS05A, __A01_1__scaler_s5__FS_n, F05A_n, __A01_1__F05A, F05B_n, __A01_1__F05B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1129(CHAT01, RCHAT_n, __A01_1__scaler_s6__FS_n, CHAT02, RCHAT_n, __A01_1__scaler_s7__FS_n, GND, RCHAT_n, __A01_1__scaler_s8__FS_n, CHAT03, RCHAT_n, __A01_1__scaler_s9__FS_n, CHAT04, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1130(CHAT05, RCHAT_n, __A01_1__scaler_s10__FS_n, CHAT06, RCHAT_n, __A01_1__scaler_s11__FS_n, GND, RCHAT_n, __A01_1__scaler_s12__FS_n, CHAT07, RCHAT_n, __A01_1__scaler_s13__FS_n, CHAT08, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1131(CHAT09, RCHAT_n, __A01_1__scaler_s14__FS_n, CHAT10, RCHAT_n, __A01_1__scaler_s15__FS_n, GND, RCHAT_n, __A01_1__scaler_s16__FS_n, CHAT11, RCHAT_n, __A01_1__scaler_s17__FS_n, CHAT12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1132(F18A, __A01_2__scaler_s18__FS_n, net_U1132_Pad3, F18B, net_U1132_Pad12, __A01_2__FS18, GND, net_U1132_Pad3, __A01_2__FS18, __A01_2__scaler_s18__FS_n, __A01_2__scaler_s18__FS_n, net_U1132_Pad12, __A01_2__FS18, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1133(F18A, F17A, net_U1132_Pad3, F17A, F18B, net_U1132_Pad12, GND, net_U1133_Pad8, __A01_2__F19A, F18A, net_U1133_Pad11, net_U1132_Pad3, net_U1132_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1134(__A01_2__F19A, __A01_2__scaler_s19__FS_n, net_U1133_Pad8, __A01_2__F19B, net_U1133_Pad11, __A01_2__FS19, GND, net_U1133_Pad8, __A01_2__FS19, __A01_2__scaler_s19__FS_n, __A01_2__scaler_s19__FS_n, net_U1133_Pad11, __A01_2__FS19, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1135(net_U1133_Pad8, F18A, __A01_2__F20A, __A01_2__F19A, net_U1135_Pad5, net_U1135_Pad6, GND, net_U1135_Pad5, net_U1135_Pad6, __A01_2__F19A, __A01_2__F20B, net_U1133_Pad11, __A01_2__F19B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1136(__A01_2__F20A, __A01_2__scaler_s20__FS_n, net_U1135_Pad6, __A01_2__F20B, net_U1135_Pad5, __A01_2__FS20, GND, net_U1135_Pad6, __A01_2__FS20, __A01_2__scaler_s20__FS_n, __A01_2__scaler_s20__FS_n, net_U1135_Pad5, __A01_2__FS20, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1137(__A01_2__F21A, __A01_2__scaler_s21__FS_n, net_U1137_Pad3, __A01_2__F21B, net_U1137_Pad12, __A01_2__FS21, GND, net_U1137_Pad3, __A01_2__FS21, __A01_2__scaler_s21__FS_n, __A01_2__scaler_s21__FS_n, net_U1137_Pad12, __A01_2__FS21, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1138(__A01_2__F21A, __A01_2__F20A, net_U1137_Pad3, __A01_2__F20A, __A01_2__F21B, net_U1137_Pad12, GND, net_U1138_Pad8, __A01_2__F22A, __A01_2__F21A, net_U1138_Pad11, net_U1137_Pad3, net_U1137_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1139(__A01_2__F22A, __A01_2__scaler_s22__FS_n, net_U1138_Pad8, __A01_2__F22B, net_U1138_Pad11, __A01_2__FS22, GND, net_U1138_Pad8, __A01_2__FS22, __A01_2__scaler_s22__FS_n, __A01_2__scaler_s22__FS_n, net_U1138_Pad11, __A01_2__FS22, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1140(net_U1138_Pad8, __A01_2__F21A, __A01_2__F23A, __A01_2__F22A, net_U1140_Pad5, net_U1140_Pad6, GND, net_U1140_Pad5, net_U1140_Pad6, __A01_2__F22A, __A01_2__F23B, net_U1138_Pad11, __A01_2__F22B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1141(__A01_2__F23A, __A01_2__scaler_s23__FS_n, net_U1140_Pad6, __A01_2__F23B, net_U1140_Pad5, __A01_2__FS23, GND, net_U1140_Pad6, __A01_2__FS23, __A01_2__scaler_s23__FS_n, __A01_2__scaler_s23__FS_n, net_U1140_Pad5, __A01_2__FS23, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1142(__A01_2__F24A, __A01_2__scaler_s24__FS_n, net_U1142_Pad3, __A01_2__F24B, net_U1142_Pad12, __A01_2__FS24, GND, net_U1142_Pad3, __A01_2__FS24, __A01_2__scaler_s24__FS_n, __A01_2__scaler_s24__FS_n, net_U1142_Pad12, __A01_2__FS24, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1143(__A01_2__F24A, __A01_2__F23A, net_U1142_Pad3, __A01_2__F23A, __A01_2__F24B, net_U1142_Pad12, GND, net_U1143_Pad8, __A01_2__F25A, __A01_2__F24A, net_U1143_Pad11, net_U1142_Pad3, net_U1142_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1144(__A01_2__F25A, __A01_2__scaler_s25__FS_n, net_U1143_Pad8, __A01_2__F25B, net_U1143_Pad11, __A01_2__FS25, GND, net_U1143_Pad8, __A01_2__FS25, __A01_2__scaler_s25__FS_n, __A01_2__scaler_s25__FS_n, net_U1143_Pad11, __A01_2__FS25, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1145(net_U1143_Pad8, __A01_2__F24A, __A01_2__F26A, __A01_2__F25A, net_U1145_Pad5, net_U1145_Pad6, GND, net_U1145_Pad5, net_U1145_Pad6, __A01_2__F25A, __A01_2__F26B, net_U1143_Pad11, __A01_2__F25B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1146(__A01_2__F26A, __A01_2__scaler_s26__FS_n, net_U1145_Pad6, __A01_2__F26B, net_U1145_Pad5, __A01_2__FS26, GND, net_U1145_Pad6, __A01_2__FS26, __A01_2__scaler_s26__FS_n, __A01_2__scaler_s26__FS_n, net_U1145_Pad5, __A01_2__FS26, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1147(__A01_2__F27A, __A01_2__scaler_s27__FS_n, net_U1147_Pad3, __A01_2__F27B, net_U1147_Pad12, __A01_2__FS27, GND, net_U1147_Pad3, __A01_2__FS27, __A01_2__scaler_s27__FS_n, __A01_2__scaler_s27__FS_n, net_U1147_Pad12, __A01_2__FS27, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1148(__A01_2__F27A, __A01_2__F26A, net_U1147_Pad3, __A01_2__F26A, __A01_2__F27B, net_U1147_Pad12, GND, net_U1148_Pad8, __A01_2__F28A, __A01_2__F27A, net_U1148_Pad11, net_U1147_Pad3, net_U1147_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1149(__A01_2__F28A, __A01_2__scaler_s28__FS_n, net_U1148_Pad8, __A01_2__F28B, net_U1148_Pad11, __A01_2__FS28, GND, net_U1148_Pad8, __A01_2__FS28, __A01_2__scaler_s28__FS_n, __A01_2__scaler_s28__FS_n, net_U1148_Pad11, __A01_2__FS28, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1150(net_U1148_Pad8, __A01_2__F27A, __A01_2__F29A, __A01_2__F28A, net_U1150_Pad5, net_U1150_Pad6, GND, net_U1150_Pad5, net_U1150_Pad6, __A01_2__F28A, __A01_2__F29B, net_U1148_Pad11, __A01_2__F28B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1151(__A01_2__F29A, __A01_2__scaler_s29__FS_n, net_U1150_Pad6, __A01_2__F29B, net_U1150_Pad5, __A01_2__FS29, GND, net_U1150_Pad6, __A01_2__FS29, __A01_2__scaler_s29__FS_n, __A01_2__scaler_s29__FS_n, net_U1150_Pad5, __A01_2__FS29, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1152(__A01_2__F30A, __A01_2__scaler_s30__FS_n, net_U1152_Pad3, __A01_2__F30B, net_U1152_Pad12, __A01_2__FS30, GND, net_U1152_Pad3, __A01_2__FS30, __A01_2__scaler_s30__FS_n, __A01_2__scaler_s30__FS_n, net_U1152_Pad12, __A01_2__FS30, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1153(__A01_2__F30A, __A01_2__F29A, net_U1152_Pad3, __A01_2__F29A, __A01_2__F30B, net_U1152_Pad12, GND, net_U1153_Pad8, __A01_2__F31A, __A01_2__F30A, net_U1153_Pad11, net_U1152_Pad3, net_U1152_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1154(__A01_2__F31A, __A01_2__scaler_s31__FS_n, net_U1153_Pad8, __A01_2__F31B, net_U1153_Pad11, __A01_2__FS31, GND, net_U1153_Pad8, __A01_2__FS31, __A01_2__scaler_s31__FS_n, __A01_2__scaler_s31__FS_n, net_U1153_Pad11, __A01_2__FS31, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1155(net_U1153_Pad8, __A01_2__F30A, __A01_2__F32A, __A01_2__F31A, net_U1155_Pad5, net_U1155_Pad6, GND, net_U1155_Pad5, net_U1155_Pad6, __A01_2__F31A, __A01_2__F32B, net_U1153_Pad11, __A01_2__F31B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1156(__A01_2__F32A, __A01_2__scaler_s32__FS_n, net_U1155_Pad6, __A01_2__F32B, net_U1155_Pad5, __A01_2__FS32, GND, net_U1155_Pad6, __A01_2__FS32, __A01_2__scaler_s32__FS_n, __A01_2__scaler_s32__FS_n, net_U1155_Pad5, __A01_2__FS32, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1157(__A01_2__F33A, __A01_2__scaler_s33__FS_n, net_U1157_Pad3, __A01_2__F33B, net_U1157_Pad12, __A01_2__FS33, GND, net_U1157_Pad3, __A01_2__FS33, __A01_2__scaler_s33__FS_n, __A01_2__scaler_s33__FS_n, net_U1157_Pad12, __A01_2__FS33, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1158(__A01_2__F33A, __A01_2__F32A, net_U1157_Pad3, __A01_2__F32A, __A01_2__F33B, net_U1157_Pad12, GND,  ,  ,  ,  , net_U1157_Pad3, net_U1157_Pad12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1159(CHAT13, RCHAT_n, __A01_2__scaler_s18__FS_n, CHAT14, RCHAT_n, __A01_2__scaler_s19__FS_n, GND, RCHBT_n, __A01_2__scaler_s20__FS_n, CHBT01, RCHBT_n, __A01_2__scaler_s21__FS_n, CHBT02, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1160(CHBT03, RCHBT_n, __A01_2__scaler_s22__FS_n, CHBT04, RCHBT_n, __A01_2__scaler_s23__FS_n, GND, RCHBT_n, __A01_2__scaler_s24__FS_n, CHBT05, RCHBT_n, __A01_2__scaler_s25__FS_n, CHBT06, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1161(CHBT07, RCHBT_n, __A01_2__scaler_s26__FS_n, CHBT08, RCHBT_n, __A01_2__scaler_s27__FS_n, GND, RCHBT_n, __A01_2__scaler_s28__FS_n, CHBT09, RCHBT_n, __A01_2__scaler_s29__FS_n, CHBT10, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1162(CHBT11, RCHBT_n, __A01_2__scaler_s30__FS_n, CHBT12, RCHBT_n, __A01_2__scaler_s31__FS_n, GND, RCHBT_n, __A01_2__scaler_s32__FS_n, CHBT13, RCHBT_n, __A01_2__scaler_s33__FS_n, CHBT14, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U1163(F07B, F07B_n, F10A, F10A_n, F09B, F09B_n, GND, FS07_n, __A01_1__FS07, FS07A, FS07_n, FS05_n, FS05, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U1164(FS09, FS09_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
endmodule