`timescale 1ns/1ps
`default_nettype none

module sq_register(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, T01_n, T02, T12_n, PHS2_n, RT_n, CT_n, WT_n, WL16_n, WL14_n, WL13_n, WL12_n, WL11_n, WL10_n, INKL, INHPLS, RELPLS, RUPTOR_n, RPTSET, KRPT, ST0_n, ST1_n, STD2, ST3_n, BR2_n, BR1B2B, RXOR0, EXT, EXTPLS, NISQ, NISQ_n, n5XP4, A15_n, A16_n, MTCSAI, MNHRPT, NISQL_n, RBSQ, SQ0_n, SQ1_n, SQ2_n, QC0_n, QC1_n, QC2_n, QC3_n, SQR12_n, SQR10, SQR10_n, SQEXT, SQEXT_n, EXST0_n, EXST1_n, FUTEXT, IIP, IIP_n, STRTFC, AD0, ADS0, AUG0_n, CCS0, CCS0_n, DAS0, DAS0_n, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DXCH0, GOJ1, GOJ1_n, INCR0, MASK0, MASK0_n, MP0, MP0_n, MP1, MP1_n, MP3, MP3_n, MP3A, MSU0, MSU0_n, NDX0_n, NDXX1_n, QXCH0_n, RSM3, RSM3_n, SU0, TC0, TC0_n, TCF0, TCSAJ3, TCSAJ3_n, TS0, TS0_n, IC1, IC2, IC2_n, IC3, IC4, IC5, IC5_n, IC6, IC7, IC8_n, IC9, IC10, IC10_n, IC11, IC11_n, IC12, IC12_n, IC13, IC14, IC15, IC15_n, IC16, IC16_n, IC17, MSQ16, MSQ14, MSQ13, MSQ12, MSQ11, MSQ10, MSQEXT, MINHL, MIIP, MTCSA_n);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire A15_n;
    input wire A16_n;
    output wire AD0;
    output wire ADS0;
    output wire AUG0_n;
    input wire BR1B2B;
    input wire BR2_n;
    output wire CCS0;
    output wire CCS0_n;
    input wire CT_n;
    output wire DAS0;
    output wire DAS0_n;
    output wire DAS1;
    output wire DAS1_n;
    output wire DCA0;
    output wire DCS0;
    output wire DIM0_n;
    output wire DXCH0;
    output wire EXST0_n;
    output wire EXST1_n;
    input wire EXT;
    input wire EXTPLS;
    output wire FUTEXT;
    output wire GOJ1;
    output wire GOJ1_n;
    input wire GOJAM;
    output wire IC1;
    output wire IC10;
    output wire IC10_n;
    output wire IC11;
    output wire IC11_n;
    output wire IC12;
    output wire IC12_n;
    output wire IC13;
    output wire IC14;
    output wire IC15;
    output wire IC15_n;
    output wire IC16;
    output wire IC16_n;
    output wire IC17;
    output wire IC2;
    output wire IC2_n;
    output wire IC3;
    output wire IC4;
    output wire IC5;
    output wire IC5_n;
    output wire IC6;
    output wire IC7;
    output wire IC8_n;
    output wire IC9;
    output wire IIP;
    output wire IIP_n;
    output wire INCR0;
    input wire INHPLS;
    input wire INKL;
    input wire KRPT;
    output wire MASK0;
    output wire MASK0_n;
    output wire MIIP; //FPGA#wand
    output wire MINHL; //FPGA#wand
    input wire MNHRPT;
    output wire MP0;
    output wire MP0_n;
    output wire MP1;
    output wire MP1_n;
    output wire MP3;
    output wire MP3A;
    output wire MP3_n;
    output wire MSQ10; //FPGA#wand
    output wire MSQ11; //FPGA#wand
    output wire MSQ12; //FPGA#wand
    output wire MSQ13; //FPGA#wand
    output wire MSQ14; //FPGA#wand
    output wire MSQ16; //FPGA#wand
    output wire MSQEXT; //FPGA#wand
    output wire MSU0;
    output wire MSU0_n;
    input wire MTCSAI;
    output wire MTCSA_n; //FPGA#wand
    output wire NDX0_n;
    output wire NDXX1_n;
    input wire NISQ;
    output wire NISQL_n;
    input wire NISQ_n;
    input wire PHS2_n;
    output wire QC0_n;
    output wire QC1_n;
    output wire QC2_n;
    output wire QC3_n;
    output wire QXCH0_n;
    output wire RBSQ;
    input wire RELPLS;
    inout wire RPTSET; //FPGA#wand
    output wire RSM3;
    output wire RSM3_n;
    input wire RT_n;
    input wire RUPTOR_n;
    input wire RXOR0;
    output wire SQ0_n;
    output wire SQ1_n;
    output wire SQ2_n;
    output wire SQEXT;
    output wire SQEXT_n;
    output wire SQR10;
    output wire SQR10_n;
    output wire SQR12_n;
    input wire ST0_n;
    input wire ST1_n;
    input wire ST3_n;
    input wire STD2;
    output wire STRTFC;
    output wire SU0;
    input wire T01_n;
    input wire T02;
    input wire T12_n;
    output wire TC0;
    output wire TC0_n;
    output wire TCF0;
    output wire TCSAJ3;
    output wire TCSAJ3_n;
    output wire TS0;
    output wire TS0_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL16_n;
    input wire WT_n;
    wire __A03_1__CSQG;
    wire __A03_1__INHINT;
    wire __A03_1__INKBT1;
    wire __A03_1__NISQL;
    wire __A03_1__OVNHRP;
    wire __A03_1__QC0;
    wire __A03_1__RPTFRC;
    wire __A03_1__SQ3_n;
    wire __A03_1__SQ4_n;
    wire __A03_1__SQ5_n;
    wire __A03_1__SQ6_n;
    wire __A03_1__SQ7_n;
    wire __A03_1__SQR11;
    wire __A03_1__SQR12;
    wire __A03_1__SQR13;
    wire __A03_1__SQR14;
    wire __A03_1__SQR16;
    wire __A03_1__WSQG_n;
    wire __A03_1__wsqg;
    wire __A03_2__AUG0;
    wire __A03_2__BMF0;
    wire __A03_2__BMF0_n;
    wire __A03_2__BZF0;
    wire __A03_2__BZF0_n;
    wire __A03_2__DIM0;
    wire __A03_2__IC13_n; //FPGA#wand
    wire __A03_2__IC3_n;
    wire __A03_2__IC4_n;
    wire __A03_2__IC9_n;
    wire __A03_2__LXCH0;
    wire __A03_2__NDX0;
    wire __A03_2__NDXX1;
    wire __A03_2__NEXST0;
    wire __A03_2__NEXST0_n;
    wire __A03_2__QXCH0;
    wire __A03_2__SQ5QC0_n;
    wire __A03_NET_163;
    wire __A03_NET_164;
    wire __A03_NET_165;
    wire __A03_NET_166;
    wire __A03_NET_167;
    wire __A03_NET_168;
    wire __A03_NET_169;
    wire __A03_NET_170;
    wire __A03_NET_171;
    wire __A03_NET_172;
    wire __A03_NET_173;
    wire __A03_NET_174;
    wire __A03_NET_175;
    wire __A03_NET_176;
    wire __A03_NET_177;
    wire __A03_NET_178;
    wire __A03_NET_179;
    wire __A03_NET_180;
    wire __A03_NET_181;
    wire __A03_NET_182;
    wire __A03_NET_183;
    wire __A03_NET_184;
    wire __A03_NET_185;
    wire __A03_NET_186;
    wire __A03_NET_187;
    wire __A03_NET_188;
    wire __A03_NET_189;
    wire __A03_NET_190;
    wire __A03_NET_191;
    wire __A03_NET_192;
    wire __A03_NET_193;
    wire __A03_NET_194;
    wire __A03_NET_196;
    wire __A03_NET_197;
    wire __A03_NET_198;
    wire __A03_NET_199;
    wire __A03_NET_200;
    wire __A03_NET_201;
    wire __A03_NET_202;
    wire __A03_NET_203;
    wire __A03_NET_204;
    wire __A03_NET_205;
    wire __A03_NET_206;
    wire __A03_NET_207;
    wire __A03_NET_208;
    wire __A03_NET_209;
    wire __A03_NET_211;
    wire __A03_NET_213;
    wire __A03_NET_214;
    wire __A03_NET_215;
    wire __A03_NET_216;
    wire __A03_NET_217;
    wire __A03_NET_218;
    wire __A03_NET_219;
    wire __A03_NET_220;
    wire __A03_NET_221;
    wire __A03_NET_223;
    wire __A03_NET_224;
    wire __A03_NET_225;
    wire __A03_NET_226;
    wire __A03_NET_227;
    wire __A03_NET_228;
    wire __A03_NET_231;
    wire __A03_NET_232;
    wire __A03_NET_234;
    wire __A03_NET_235;
    wire __A03_NET_236;
    wire __A03_NET_237;
    wire __A03_NET_238;
    wire __A03_NET_239;
    wire __A03_NET_240;
    wire __A03_NET_242;
    input wire n5XP4;

    pullup R3001(RPTSET);
    pullup R3002(__A03_2__IC13_n);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U3001(__A03_NET_211, NISQ, __A03_1__NISQL, __A03_NET_213, STRTFC, __A03_NET_220, GND, RT_n, __A03_NET_209, RBSQ, __A03_NET_209, WT_n, __A03_1__wsqg, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3002(__A03_NET_211, __A03_1__INKBT1, T12_n, __A03_NET_211, __A03_1__RPTFRC, __A03_NET_220, GND, __A03_1__CSQG, T12_n, CT_n, __A03_NET_213, __A03_1__NISQL, STRTFC, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U3003(__A03_1__NISQL, NISQL_n, __A03_NET_220, __A03_NET_209, __A03_1__wsqg, __A03_1__WSQG_n, GND, STRTFC, __A03_NET_217, SQEXT, __A03_NET_216, SQEXT_n, __A03_NET_221, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U3004(__A03_NET_165, WL16_n, __A03_1__WSQG_n, __A03_NET_166, WL14_n, __A03_1__WSQG_n, GND, WL13_n, __A03_1__WSQG_n, __A03_NET_167, __A03_NET_190, __A03_NET_187, __A03_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3005(__A03_NET_217, GOJAM, MTCSAI, __A03_NET_218, NISQL_n, T12_n, GND, STRTFC, __A03_NET_218, __A03_NET_219, __A03_NET_219, __A03_NET_182, __A03_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U3006(EXTPLS, EXT, __A03_NET_182, __A03_1__INKBT1, STRTFC, FUTEXT, GND, __A03_NET_216, __A03_1__RPTFRC, __A03_NET_215, __A03_NET_221, __A03_NET_182, FUTEXT, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U3007(__A03_NET_214, __A03_NET_219, FUTEXT, __A03_NET_221, __A03_NET_216, __A03_NET_214, GND, INHPLS, __A03_1__INHINT, __A03_NET_180, KRPT, IIP, IIP_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3009(__A03_NET_180, RELPLS, IIP_n, GOJAM, n5XP4, IIP, GND, __A03_NET_178, FUTEXT, NISQL_n, T12_n, __A03_1__INHINT, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3010(PHS2_n, RUPTOR_n, __A03_1__OVNHRP, __A03_1__INHINT, IIP, __A03_NET_177, GND, __A03_NET_183, __A03_NET_181, STRTFC, T02, __A03_NET_179, MNHRPT, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U3011(__A03_NET_178, RPTSET, __A03_NET_179, RPTSET, __A03_NET_177, RPTSET, GND, __A03_2__IC13_n, __A03_NET_238, __A03_2__IC13_n, __A03_NET_239,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U3012(__A03_NET_181, RPTSET, __A03_NET_183, __A03_NET_192, __A03_NET_165, __A03_1__SQR16, GND, __A03_NET_166, __A03_1__SQR14, __A03_NET_193, __A03_NET_167, __A03_1__SQR13, __A03_NET_194, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3013(__A03_NET_192, __A03_1__RPTFRC, __A03_NET_193, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR14, GND, __A03_1__SQR13, __A03_NET_194, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR16, __A03_1__CSQG, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U3014(__A03_NET_163, __A03_NET_192, INKL, __A03_NET_164, INKL, __A03_1__SQR16, GND, __A03_NET_184, __A03_1__OVNHRP, __A03_NET_189, __A03_NET_185, NISQ_n, __A03_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U3015(__A03_NET_198, __A03_NET_168, __A03_NET_194, __A03_NET_168, __A03_NET_175, __A03_NET_169, GND, __A03_NET_170, __A03_NET_198, __A03_NET_193, __A03_NET_175, __A03_NET_176, __A03_NET_175, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3016(__A03_NET_194, __A03_NET_193, __A03_NET_198, __A03_NET_168, __A03_NET_199, __A03_NET_172, GND, __A03_NET_204, __A03_NET_194, __A03_NET_168, __A03_NET_199, __A03_NET_171, __A03_NET_175, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U3017(__A03_NET_198, __A03_NET_199, __A03_NET_194, __A03_NET_193, __A03_NET_199, __A03_NET_174, GND, __A03_NET_205, __A03_1__RPTFRC, __A03_NET_200, __A03_1__SQR12, __A03_NET_173, __A03_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3018(__A03_NET_169, SQ1_n, __A03_NET_170, SQ2_n, __A03_NET_171, __A03_1__SQ3_n, GND, __A03_1__SQ4_n, __A03_NET_172, __A03_1__SQ6_n, __A03_NET_173, __A03_1__SQ7_n, __A03_NET_174, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3019(__A03_NET_200, WL12_n, __A03_1__WSQG_n, __A03_NET_197, WL11_n, __A03_1__WSQG_n, GND, __A03_NET_205, __A03_1__CSQG, __A03_1__SQR12, __A03_NET_196, __A03_1__CSQG, __A03_1__SQR11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U3020(__A03_1__RPTFRC, __A03_NET_197, __A03_1__RPTFRC, __A03_NET_201, __A03_NET_202, __A03_NET_203, GND, __A03_1__INKBT1, INKL, T01_n, STD2, __A03_NET_196, __A03_1__SQR11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3021(A16_n, __A03_NET_188, A15_n, __A03_NET_186,  ,  , GND, SQR12_n, __A03_1__SQR12, __A03_1__RPTFRC, __A03_NET_181, __A03_1__SQ5_n, __A03_NET_204, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3022(__A03_1__QC0, __A03_1__SQR11, __A03_1__SQR12, __A03_NET_206, __A03_NET_196, __A03_1__SQR12, GND, __A03_1__SQR11, __A03_NET_205, __A03_NET_207, __A03_NET_205, __A03_NET_196, __A03_NET_208, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3023(__A03_1__QC0, QC0_n, __A03_NET_206, QC1_n, __A03_NET_207, QC2_n, GND, QC3_n, __A03_NET_208, SQR10, __A03_NET_203, SQR10_n, __A03_NET_202, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3024(__A03_NET_201, WL10_n, __A03_1__WSQG_n, __A03_NET_202, __A03_NET_203, __A03_1__CSQG, GND, __A03_NET_188, A15_n, __A03_NET_190, A16_n, __A03_NET_186, __A03_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3025(__A03_NET_163, __A03_NET_199, __A03_NET_164, __A03_NET_175, __A03_NET_193, __A03_NET_168, GND, __A03_NET_198, __A03_NET_194, SQ0_n, __A03_NET_176, MP3A, MP3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3026(__A03_NET_235, __A03_1__SQ5_n, QC0_n, __A03_NET_236, __A03_1__SQ5_n, SQEXT_n, GND, __A03_NET_235, __A03_NET_236, __A03_NET_242, __A03_NET_242, ST0_n, IC1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U3027(__A03_NET_235, __A03_2__SQ5QC0_n, IC2, IC2_n, __A03_NET_228, EXST1_n, GND, TC0_n, TC0, IC3, __A03_2__IC3_n, __A03_2__NEXST0_n, __A03_2__NEXST0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3028(IC2, __A03_NET_242, ST1_n, __A03_NET_237, SQEXT_n, __A03_1__QC0, GND, SQEXT_n, ST1_n, __A03_NET_228, __A03_NET_228, __A03_2__NEXST0, __A03_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3029(__A03_NET_237, __A03_1__SQ6_n, SQ1_n, __A03_2__NEXST0_n, __A03_1__QC0, TCF0, GND, __A03_2__IC3_n, TC0, STD2, TCF0, IC11, ST0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3030(IC6, __A03_NET_234, __A03_1__SQ3_n, IC7, __A03_NET_234, __A03_1__SQ4_n, GND, SQ0_n, __A03_2__NEXST0_n, TC0, SQEXT, ST0_n, __A03_2__NEXST0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3031(DCS0, __A03_1__SQ4_n, EXST0_n, DCA0, EXST0_n, __A03_1__SQ3_n, GND, DCS0, DCA0, __A03_2__IC4_n, QC1_n, ST1_n, __A03_NET_240, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3032(IC7, IC6, IC1, DCS0, DCA0, __A03_NET_239, GND, IC5, __A03_NET_231, __A03_1__SQ5_n, SQEXT, __A03_NET_238, IC11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3033(__A03_2__IC4_n, IC4, __A03_2__IC13_n, IC13, IC5, IC5_n, GND, IC9, __A03_2__IC9_n, QXCH0_n, __A03_2__QXCH0, EXST0_n, __A03_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3034(__A03_NET_232, QC3_n, ST0_n, __A03_NET_231, __A03_NET_240, __A03_NET_232, GND, __A03_2__LXCH0, DXCH0, IC8_n, ST0_n, SQEXT_n, __A03_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3035(__A03_2__NEXST0_n, QC1_n, SQ2_n, QC1_n, EXST0_n, __A03_2__QXCH0, GND, TS0, __A03_1__SQ5_n, QC2_n, __A03_2__NEXST0_n, __A03_2__LXCH0, SQ2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U3036(__A03_2__IC9_n, IC5, TS0, __A03_2__QXCH0, __A03_2__LXCH0,  , GND,  , SQ2_n, QC0_n, SQEXT, ST1_n, __A03_NET_224, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3037(TS0, TS0_n, IC10_n, IC10, DAS0, DAS0_n, GND, __A03_2__BZF0_n, __A03_2__BZF0, __A03_2__BMF0_n, __A03_2__BMF0, IC16, IC16_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3038(__A03_1__SQ5_n, __A03_2__NEXST0_n, SQ2_n, __A03_2__NEXST0_n, QC0_n, DAS0, GND, IC10_n, IC4, DXCH0, DAS0, DXCH0, QC1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3039(SQ1_n, __A03_1__QC0, EXST0_n, __A03_1__QC0, __A03_1__SQ6_n, __A03_2__BMF0, GND, CCS0, SQ1_n, QC0_n, __A03_2__NEXST0_n, __A03_2__BZF0, EXST0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3040(IC15_n, __A03_2__BMF0, __A03_2__BZF0, __A03_NET_226, __A03_2__BZF0_n, BR2_n, GND, __A03_2__BMF0_n, BR1B2B, __A03_NET_225, __A03_NET_226, __A03_NET_225, IC16_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U3041(IC17, IC16, IC15_n, DAS1_n, __A03_NET_224, ADS0, GND, CCS0, MSU0, IC12_n, __A03_1__SQ7_n, __A03_2__NEXST0_n, MASK0, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3042(IC15_n, IC15, CCS0, CCS0_n, DAS1_n, DAS1, GND, IC12, IC12_n, MSU0_n, MSU0, AUG0_n, __A03_2__AUG0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U3043(SQ2_n, QC3_n, QC2_n, SQ2_n, __A03_2__NEXST0_n, INCR0, GND, MSU0, SQ2_n, EXST0_n, QC0_n, ADS0, __A03_2__NEXST0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3044(SQ2_n, EXST0_n, SQ2_n, EXST0_n, QC3_n, __A03_2__DIM0, GND, MP3, ST3_n, __A03_1__SQ7_n, SQEXT_n, __A03_2__AUG0, QC2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U3045(__A03_2__DIM0, DIM0_n, MP3, MP3_n, MP1, MP1_n, GND, MP0_n, MP0, TCSAJ3_n, TCSAJ3, RSM3_n, RSM3, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3046(ST1_n, __A03_1__SQ7_n, ST0_n, __A03_1__SQ7_n, SQEXT_n, MP0, GND, TCSAJ3, SQ0_n, SQEXT, ST3_n, MP1, SQEXT_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3047(ST3_n, __A03_2__SQ5QC0_n, __A03_1__SQ6_n, EXST0_n, QC0_n, SU0, GND, __A03_NET_227, MP0, MASK0, RXOR0, RSM3, SQEXT, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3048(MASK0, MASK0_n, __A03_NET_227, IC14, __A03_2__NDX0, NDX0_n, GND, NDXX1_n, __A03_2__NDXX1, GOJ1_n, GOJ1, IC11_n, IC11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3049(AD0, __A03_2__NEXST0_n, __A03_1__SQ6_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3050(__A03_2__NEXST0_n, __A03_1__SQ5_n, SQEXT_n, __A03_1__SQ5_n, ST1_n, __A03_2__NDXX1, GND, GOJ1, SQEXT, ST1_n, SQ0_n, __A03_2__NDX0, QC0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3052(__A03_NET_189, __A03_NET_191, __A03_NET_190, __A03_NET_187, NISQ_n, __A03_NET_191, GND,  ,  ,  ,  , __A03_1__OVNHRP, MP3, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U3053(__A03_NET_203, MSQ10, __A03_NET_180, MINHL, IIP_n, MIIP, GND, MTCSA_n, TCSAJ3,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8
    U74LVC06 U3054(__A03_NET_216, MSQEXT, __A03_NET_192, MSQ16, __A03_NET_193, MSQ14, GND, MSQ13, __A03_NET_194, MSQ12, __A03_NET_205, MSQ11, __A03_NET_196, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
endmodule