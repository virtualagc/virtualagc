`timescale 1ns/1ps
`default_nettype none

module fixed_erasable_memory(SIM_RST, SIM_CLK, p4VSW, GND, ROPER, ROPES, ROPET, HIMOD, LOMOD, STR14, STR58, STR912, STR19, STR210, STR311, STR412, SETAB, SETCD, RESETA, RESETB, RESETC, RESETD, CLROPE, IL07, IL06, IL05, IL04, IL03, IL02, IL01, SBF, XB7E, XB1E, XB2E, XB3E, XB4E, XB5E, XB6E, XT7E, XT1E, XT2E, XT3E, XT4E, XT5E, XT6E, YB3E, YB1E, YB2E, YT7E, YT1E, YT2E, YT3E, YT4E, YT5E, YT6E, GEMP, GEM01, GEM02, GEM03, GEM04, GEM05, GEM06, GEM07, GEM08, GEM09, GEM10, GEM11, GEM12, GEM13, GEM14, GEM16, SETEK, RSTKX_n, RSTKY_n, SBE, REX, REY, WEX, WEY, ZID, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08, SA09, SA10, SA11, SA12, SA13, SA14, SAP, SA16);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire CLROPE;
    input wire GEM01;
    input wire GEM02;
    input wire GEM03;
    input wire GEM04;
    input wire GEM05;
    input wire GEM06;
    input wire GEM07;
    input wire GEM08;
    input wire GEM09;
    input wire GEM10;
    input wire GEM11;
    input wire GEM12;
    input wire GEM13;
    input wire GEM14;
    input wire GEM16;
    input wire GEMP;
    input wire HIMOD;
    input wire IL01;
    input wire IL02;
    input wire IL03;
    input wire IL04;
    input wire IL05;
    input wire IL06;
    input wire IL07;
    input wire LOMOD;
    input wire RESETA;
    input wire RESETB;
    input wire RESETC;
    input wire RESETD;
    input wire REX;
    input wire REY;
    input wire ROPER;
    input wire ROPES;
    input wire ROPET;
    input wire RSTKX_n;
    input wire RSTKY_n;
    output wire SA01; //FPGA#wor
    output wire SA02; //FPGA#wor
    output wire SA03; //FPGA#wor
    output wire SA04; //FPGA#wor
    output wire SA05; //FPGA#wor
    output wire SA06; //FPGA#wor
    output wire SA07; //FPGA#wor
    output wire SA08; //FPGA#wor
    output wire SA09; //FPGA#wor
    output wire SA10; //FPGA#wor
    output wire SA11; //FPGA#wor
    output wire SA12; //FPGA#wor
    output wire SA13; //FPGA#wor
    output wire SA14; //FPGA#wor
    output wire SA16; //FPGA#wor
    output wire SAP; //FPGA#wor
    input wire SBE;
    input wire SBF;
    input wire SETAB;
    input wire SETCD;
    input wire SETEK;
    input wire STR14;
    input wire STR19;
    input wire STR210;
    input wire STR311;
    input wire STR412;
    input wire STR58;
    input wire STR912;
    input wire WEX;
    input wire WEY;
    input wire XB1E;
    input wire XB2E;
    input wire XB3E;
    input wire XB4E;
    input wire XB5E;
    input wire XB6E;
    input wire XB7E;
    input wire XT1E;
    input wire XT2E;
    input wire XT3E;
    input wire XT4E;
    input wire XT5E;
    input wire XT6E;
    input wire XT7E;
    input wire YB1E;
    input wire YB2E;
    input wire YB3E;
    input wire YT1E;
    input wire YT2E;
    input wire YT3E;
    input wire YT4E;
    input wire YT5E;
    input wire YT6E;
    input wire YT7E;
    input wire ZID;
    wire __B01_1__CQA;
    wire __B01_1__CQB;
    wire __B01_1__CQC;
    wire __B01_1__FADDR1;
    wire __B01_1__FADDR10;
    wire __B01_1__FADDR11;
    wire __B01_1__FADDR12;
    wire __B01_1__FADDR13;
    wire __B01_1__FADDR14;
    wire __B01_1__FADDR15;
    wire __B01_1__FADDR16;
    wire __B01_1__FADDR2;
    wire __B01_1__FADDR3;
    wire __B01_1__FADDR4;
    wire __B01_1__FADDR5;
    wire __B01_1__FADDR6;
    wire __B01_1__FADDR7;
    wire __B01_1__FADDR8;
    wire __B01_1__FADDR9;
    wire __B01_1__NOROPE;
    wire __B01_1__QUARTERA;
    wire __B01_1__QUARTERB;
    wire __B01_1__QUARTERC;
    wire __B01_2__EDESTROY;
    wire __B01_2__ES01_n;
    wire __B01_2__ES02_n;
    wire __B01_2__ES03_n;
    wire __B01_2__ES04_n;
    wire __B01_2__ES05_n;
    wire __B01_2__ES06_n;
    wire __B01_2__ES07_n;
    wire __B01_2__ES08_n;
    wire __B01_2__ES09_n;
    wire __B01_2__ES10_n;
    wire __B01_2__ES11_n;
    wire __B01_2__RADDR1;
    wire __B01_2__RADDR10;
    wire __B01_2__RADDR11;
    wire __B01_2__RADDR2;
    wire __B01_2__RADDR3;
    wire __B01_2__RADDR4;
    wire __B01_2__RADDR5;
    wire __B01_2__RADDR6;
    wire __B01_2__RADDR7;
    wire __B01_2__RADDR8;
    wire __B01_2__RADDR9;
    wire __B01_2__RESETK;
    wire net_U31001_Pad26;
    wire net_U31001_Pad28;
    wire net_U31002_Pad10;
    wire net_U31002_Pad12;
    wire net_U31002_Pad2;
    wire net_U31002_Pad4;
    wire net_U31002_Pad6;
    wire net_U31002_Pad8;
    wire net_U31003_Pad4;
    wire net_U31003_Pad5;
    wire net_U31004_Pad6;
    wire net_U31004_Pad8;
    wire net_U31005_Pad1;
    wire net_U31005_Pad10;
    wire net_U31005_Pad13;
    wire net_U31005_Pad4;
    wire net_U31006_Pad10;
    wire net_U31006_Pad11;
    wire net_U31006_Pad12;
    wire net_U31006_Pad9;
    wire net_U31010_Pad11;
    wire net_U31010_Pad12;
    wire net_U31010_Pad13;
    wire net_U31010_Pad4;
    wire net_U31012_Pad10;
    wire net_U31012_Pad11;
    wire net_U31012_Pad12;
    wire net_U31012_Pad13;
    wire net_U31012_Pad3;
    wire net_U31014_Pad1;
    wire net_U31014_Pad12;
    wire net_U31014_Pad13;
    wire net_U31014_Pad3;
    wire net_U31014_Pad4;
    wire net_U31015_Pad10;
    wire net_U31015_Pad11;
    wire net_U31015_Pad12;
    wire net_U31015_Pad2;
    wire net_U31015_Pad4;
    wire net_U31015_Pad5;
    wire net_U31015_Pad6;
    wire net_U31016_Pad11;
    wire net_U31016_Pad12;
    wire net_U31016_Pad6;
    wire net_U31016_Pad8;
    wire net_U31017_Pad1;
    wire net_U31017_Pad10;
    wire net_U31017_Pad8;
    wire net_U31025_Pad17;
    wire net_U31025_Pad41;
    wire net_U31026_Pad1;
    wire net_U31026_Pad10;
    wire net_U31026_Pad2;
    wire net_U31026_Pad3;
    wire net_U31026_Pad4;
    wire net_U31026_Pad6;
    wire net_U31027_Pad12;
    wire net_U31027_Pad13;
    wire net_U31027_Pad5;
    wire net_U31027_Pad6;
    wire net_U31028_Pad1;
    wire net_U31028_Pad13;
    wire net_U31028_Pad4;
    wire net_U31029_Pad1;
    wire net_U31029_Pad10;
    wire net_U31029_Pad13;
    wire net_U31030_Pad10;
    wire net_U31030_Pad4;
    wire net_U31031_Pad1;
    wire net_U31031_Pad13;
    wire net_U31031_Pad4;
    wire net_U31032_Pad1;
    wire net_U31032_Pad10;
    wire net_U31032_Pad13;
    wire net_U31033_Pad10;
    wire net_U31033_Pad4;
    wire net_U31034_Pad1;
    wire net_U31034_Pad13;
    wire net_U31034_Pad4;
    wire net_U31035_Pad1;
    wire net_U31035_Pad13;
    wire net_U31035_Pad4;
    wire net_U31035_Pad6;
    wire net_U31035_Pad9;
    wire net_U31036_Pad10;
    wire net_U31037_Pad10;
    wire net_U31037_Pad11;
    wire net_U31037_Pad12;
    wire net_U31037_Pad6;
    wire net_U31038_Pad10;
    wire net_U31038_Pad11;
    wire net_U31038_Pad12;
    wire net_U31038_Pad3;
    wire net_U31038_Pad5;
    wire net_U31038_Pad6;
    wire net_U31039_Pad10;
    wire net_U31039_Pad3;
    wire net_U31040_Pad11;

    pulldown R31001(SA01);
    pulldown R31002(SA02);
    pulldown R31003(SA03);
    pulldown R31004(SA04);
    pulldown R31005(SA05);
    pulldown R31006(SA06);
    pulldown R31007(SA07);
    pulldown R31008(SA08);
    pulldown R31009(SA09);
    pulldown R31010(SA10);
    pulldown R31011(SA11);
    pulldown R31012(SA12);
    pulldown R31013(SA13);
    pulldown R31014(SA14);
    pulldown R31015(SAP);
    pulldown R31016(SA16);
    SST39VF200A U31001(__B01_1__FADDR16, __B01_1__FADDR15, __B01_1__FADDR14, __B01_1__FADDR13, __B01_1__FADDR12, __B01_1__FADDR11, __B01_1__FADDR10, __B01_1__FADDR9,  ,  , p4VSW,  ,  ,  ,  ,  ,  , __B01_1__FADDR8, __B01_1__FADDR7, __B01_1__FADDR6, __B01_1__FADDR5, __B01_1__FADDR4, __B01_1__FADDR3, __B01_1__FADDR2, __B01_1__FADDR1, net_U31001_Pad26, GND, net_U31001_Pad28, SA01, SA09, SA02, SA10, SA03, SA11, SA04, SA12, p4VSW, SA05, SA13, SA06, SA14, SA07, SAP, SA08, SA16, GND,  , GND, SIM_RST, SIM_CLK); //FPGA#inputs:EPCS_DATA;FPGA#outputs:EPCS_CSN,EPCS_DCLK,EPCS_ASDI;FPGA#OD:29,30,31,32,33,34,35,36,38,39,40,41,42,43,44,45
    U74HC04 U31002(ROPER, net_U31002_Pad2, ROPES, net_U31002_Pad4, ROPET, net_U31002_Pad6, GND, net_U31002_Pad8, STR14, net_U31002_Pad10, STR58, net_U31002_Pad12, STR912, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31003(net_U31002_Pad6, LOMOD, ROPER, net_U31003_Pad4, net_U31003_Pad5, __B01_1__FADDR15, GND, net_U31003_Pad4, ROPES, LOMOD, STR14, __B01_1__FADDR16, STR14, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31004(ROPET, HIMOD, ROPER, LOMOD, STR14, net_U31004_Pad6, GND, net_U31004_Pad8, ROPET, LOMOD, net_U31002_Pad8, net_U31003_Pad5, STR912, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U31005(net_U31005_Pad1, net_U31002_Pad4, net_U31002_Pad12, net_U31005_Pad4, net_U31002_Pad2, HIMOD, GND, HIMOD, STR58, net_U31005_Pad10, LOMOD, net_U31002_Pad10, net_U31005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31006(__B01_1__FADDR14, net_U31005_Pad1, net_U31004_Pad6, net_U31004_Pad8, net_U31005_Pad4,  , GND,  , net_U31006_Pad9, net_U31006_Pad10, net_U31006_Pad11, net_U31006_Pad12, __B01_1__FADDR13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31007(ROPES, HIMOD, ROPES, LOMOD, STR14, net_U31006_Pad10, GND, net_U31006_Pad11, net_U31002_Pad4, HIMOD, net_U31002_Pad12, net_U31006_Pad9, STR912, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31008(net_U31002_Pad4, LOMOD, RSTKX_n, RSTKY_n, ZID, __B01_2__RESETK, GND, __B01_1__NOROPE, ROPER, ROPES, ROPET, net_U31006_Pad12, net_U31002_Pad8, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U31009(__B01_1__FADDR12, net_U31005_Pad10, net_U31005_Pad13, __B01_1__FADDR11, STR210, STR19, GND, STR19, STR311, __B01_1__FADDR10, __B01_1__QUARTERB, __B01_1__QUARTERA, __B01_1__FADDR9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31010(__B01_1__FADDR8, __B01_1__QUARTERA, __B01_1__QUARTERC, net_U31010_Pad4, net_U31010_Pad13, __B01_1__QUARTERA, GND, net_U31010_Pad4, __B01_1__CQA, __B01_1__QUARTERA, net_U31010_Pad11, net_U31010_Pad12, net_U31010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U31011(IL07, __B01_1__FADDR7, IL06, __B01_1__FADDR6, IL05, __B01_1__FADDR5, GND, __B01_1__FADDR4, IL04, __B01_1__FADDR3, IL03, __B01_1__FADDR2, IL02, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1) U31012(IL01, __B01_1__FADDR1, net_U31012_Pad3, net_U31001_Pad28, SETAB, net_U31010_Pad11, GND, net_U31010_Pad12, RESETB, net_U31012_Pad10, net_U31012_Pad11, net_U31012_Pad12, net_U31012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U31013(net_U31001_Pad26, STR19, STR210, STR311, STR412,  , GND,  , XB1E, XB3E, XB5E, XB7E, __B01_2__ES01_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31014(net_U31014_Pad1, RESETA, net_U31014_Pad3, net_U31014_Pad4, net_U31014_Pad1, net_U31012_Pad13, GND, net_U31014_Pad4, RESETA, net_U31012_Pad13, net_U31010_Pad11, net_U31014_Pad12, net_U31014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1) U31015(net_U31012_Pad12, net_U31015_Pad2, net_U31015_Pad2, net_U31015_Pad4, net_U31015_Pad5, net_U31015_Pad6, GND, net_U31015_Pad11, net_U31015_Pad6, net_U31015_Pad10, net_U31015_Pad11, net_U31015_Pad12, net_U31015_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1) U31016(net_U31015_Pad4, net_U31014_Pad3, RESETA, net_U31014_Pad12, SETCD, net_U31016_Pad6, GND, net_U31016_Pad8, RESETD, __B01_1__CQA, net_U31016_Pad11, net_U31016_Pad12, ZID, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U31017(net_U31017_Pad1, net_U31014_Pad13, __B01_1__QUARTERB, __B01_1__QUARTERB, net_U31017_Pad1, __B01_1__CQB, GND, net_U31017_Pad8, __B01_1__QUARTERC, net_U31017_Pad10, net_U31017_Pad10, __B01_1__CQC, __B01_1__QUARTERC, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U31018(net_U31017_Pad8, net_U31016_Pad6, net_U31016_Pad8, net_U31016_Pad11, CLROPE, net_U31014_Pad1, GND, YB1E, YB3E, __B01_2__ES07_n, YB2E, YB3E, __B01_2__ES08_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31019(__B01_2__ES02_n, XB2E, XB3E, XB6E, XB7E,  , GND,  , XB4E, XB5E, XB6E, XB7E, __B01_2__ES03_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31020(__B01_2__ES04_n, XT1E, XT3E, XT5E, XT7E,  , GND,  , XT2E, XT3E, XT6E, XT7E, __B01_2__ES05_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31021(__B01_2__ES06_n, XT4E, XT5E, XT6E, XT7E,  , GND,  , YT1E, YT3E, YT5E, YT7E, __B01_2__ES09_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31022(__B01_2__ES10_n, YT2E, YT3E, YT6E, YT7E,  , GND,  , YT4E, YT5E, YT6E, YT7E, __B01_2__ES11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC244 U31023(net_U31016_Pad12, GEMP, SA07, GEM01, SA06, GEM02, SA05, GEM03, SA04, GND, GEM04, SA03, GEM05, SA02, GEM06, SA01, GEM07, SAP, net_U31016_Pad12, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:3,5,7,9,12,14,16,18
    U74HC244 U31024(net_U31016_Pad12, GEM08, SA16, GEM09, SA14, GEM10, SA13, GEM11, SA12, GND, GEM12, SA11, GEM13, SA10, GEM14, SA09, GEM16, SA08, net_U31016_Pad12, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:3,5,7,9,12,14,16,18
    MR0A16A U31025(__B01_2__RADDR1, __B01_2__RADDR2, __B01_2__RADDR3, __B01_2__RADDR4, __B01_2__RADDR5, GND, SA01, SA02, SA03, SA04, p4VSW, GND, SA05, SA06, SA07, SA08, net_U31025_Pad17, __B01_2__RADDR6, __B01_2__RADDR7, __B01_2__RADDR8, __B01_2__RADDR9, __B01_2__RADDR10, __B01_2__RADDR11, GND, GND, GND, p4VSW,  , SA09, SA10, SA11, SA12, p4VSW, GND, SA13, SA14, SAP, SA16, GND, GND, net_U31025_Pad41, GND, GND, GND, SIM_RST, SIM_CLK); //FPGA#bidir:7,8,9,10,13,14,15,16,29,30,31,32,35,36,37,38;FPGA#OD:7,8,9,10,13,14,15,16,29,30,31,32,35,36,37,38
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31026(net_U31026_Pad1, net_U31026_Pad2, net_U31026_Pad3, net_U31026_Pad4, __B01_2__ES01_n, net_U31026_Pad6, GND, net_U31026_Pad4, __B01_2__RADDR1, net_U31026_Pad10, net_U31026_Pad10, __B01_2__RESETK, __B01_2__RADDR1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1) U31027(WEX, net_U31026_Pad2, WEY, net_U31026_Pad3, net_U31027_Pad5, net_U31027_Pad6, GND, net_U31025_Pad41, SBE, net_U31026_Pad6, SETEK, net_U31027_Pad12, net_U31027_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31028(net_U31028_Pad1, __B01_2__ES02_n, net_U31026_Pad6, net_U31028_Pad4, net_U31028_Pad1, __B01_2__RADDR2, GND, net_U31028_Pad4, __B01_2__RESETK, __B01_2__RADDR2, __B01_2__ES03_n, net_U31026_Pad6, net_U31028_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31029(net_U31029_Pad1, net_U31028_Pad13, __B01_2__RADDR3, __B01_2__RADDR3, net_U31029_Pad1, __B01_2__RESETK, GND, __B01_2__ES04_n, net_U31026_Pad6, net_U31029_Pad10, net_U31029_Pad10, __B01_2__RADDR4, net_U31029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31030(__B01_2__RADDR4, net_U31029_Pad13, __B01_2__RESETK, net_U31030_Pad4, __B01_2__ES05_n, net_U31026_Pad6, GND, net_U31030_Pad4, __B01_2__RADDR5, net_U31030_Pad10, net_U31030_Pad10, __B01_2__RESETK, __B01_2__RADDR5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31031(net_U31031_Pad1, __B01_2__ES06_n, net_U31026_Pad6, net_U31031_Pad4, net_U31031_Pad1, __B01_2__RADDR6, GND, net_U31031_Pad4, __B01_2__RESETK, __B01_2__RADDR6, __B01_2__ES07_n, net_U31026_Pad6, net_U31031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31032(net_U31032_Pad1, net_U31031_Pad13, __B01_2__RADDR7, __B01_2__RADDR7, net_U31032_Pad1, __B01_2__RESETK, GND, __B01_2__ES08_n, net_U31026_Pad6, net_U31032_Pad10, net_U31032_Pad10, __B01_2__RADDR8, net_U31032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31033(__B01_2__RADDR8, net_U31032_Pad13, __B01_2__RESETK, net_U31033_Pad4, __B01_2__ES09_n, net_U31026_Pad6, GND, net_U31033_Pad4, __B01_2__RADDR9, net_U31033_Pad10, net_U31033_Pad10, __B01_2__RESETK, __B01_2__RADDR9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31034(net_U31034_Pad1, __B01_2__ES10_n, net_U31026_Pad6, net_U31034_Pad4, net_U31034_Pad1, __B01_2__RADDR10, GND, net_U31034_Pad4, __B01_2__RESETK, __B01_2__RADDR10, __B01_2__ES11_n, net_U31026_Pad6, net_U31034_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31035(net_U31035_Pad1, net_U31034_Pad13, __B01_2__RADDR11, net_U31035_Pad4, CLROPE, net_U31035_Pad6, GND, net_U31027_Pad6, net_U31035_Pad9, __B01_2__EDESTROY, __B01_2__EDESTROY, net_U31027_Pad13, net_U31035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31036(net_U31027_Pad13, net_U31035_Pad13, net_U31027_Pad6, net_U31035_Pad6, RESETB, net_U31015_Pad12, GND, net_U31035_Pad6, net_U31015_Pad5, net_U31036_Pad10, net_U31036_Pad10, RESETB, net_U31015_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31037(net_U31027_Pad12, net_U31012_Pad11, net_U31035_Pad4, __B01_1__CQB, net_U31012_Pad10, net_U31037_Pad6, GND, net_U31037_Pad11, net_U31037_Pad6, net_U31037_Pad10, net_U31037_Pad11, net_U31037_Pad12, net_U31037_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31038(net_U31037_Pad12, net_U31035_Pad9, net_U31038_Pad3, __B01_1__CQC, net_U31038_Pad5, net_U31038_Pad6, GND, net_U31038_Pad11, net_U31038_Pad6, net_U31038_Pad10, net_U31038_Pad11, net_U31038_Pad12, net_U31038_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31039(net_U31038_Pad3, CLROPE, net_U31039_Pad3, net_U31039_Pad3, RESETC, net_U31038_Pad12, GND, net_U31039_Pad3, net_U31038_Pad5, net_U31039_Pad10, net_U31039_Pad10, RESETC, net_U31038_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U31040(__B01_2__RADDR11, net_U31035_Pad1, __B01_2__RESETK, net_U31027_Pad5, REX, REY, GND, net_U31026_Pad1, __B01_2__EDESTROY, net_U31025_Pad17, net_U31040_Pad11, __B01_1__NOROPE, net_U31012_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U31041(SBF, net_U31040_Pad11,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule