`timescale 1ns/1ps
`default_nettype none

module inout_iv(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, T06_n, SB0_n, SB1_n, SB2, SB2_n, F04A, F05A_n, F05B_n, F06B, FS07A, FS07_n, F07B, F09B_n, FS10, F10A_n, F10B, BR1, BR1_n, CCHG_n, CSG, POUT_n, MOUT_n, ZOUT_n, OVF_n, WOVR_n, SHINC_n, CAURST, T6ON_n, BLKUPL_n, UPL0, UPL1, XLNK0, XLNK1, GTONE, GTSET, GTSET_n, GATEX_n, GATEY_n, GATEZ_n, SIGNX, SIGNY, SIGNZ, BMGXP, BMGXM, BMGYP, BMGYM, BMGZP, BMGZM, C45R, XB3_n, XB5_n, XB6_n, XB7_n, XT3_n, CXB0_n, CXB7_n, CA2_n, CA4_n, CA5_n, CA6_n, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CCH11, CCH13, CCH14, RCH11_n, RCH13_n, RCH14_n, RCH33_n, WCH11_n, WCH13_n, WCH14_n, F5ASB0_n, F5ASB2, F5ASB2_n, F5BSB2_n, ERRST, T1P, T2P, T3P, T4P, T5P, T6P, ALTM, BMAGXP, BMAGXM, BMAGYP, BMAGYM, BMAGZP, BMAGZM, EMSD, GYROD, UPRUPT, INLNKP, INLNKM, OTLNKM, THRSTD, CCH33, CH1305, CH1306, CH1308, CH1309, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406, CH1407, CH1408, CH1409, CH1410, CH3310, CH3311, CH1109, CH1110, CH1111, CH1112);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    output wire ALTM;
    input wire BLKUPL_n;
    output wire BMAGXM;
    output wire BMAGXP;
    output wire BMAGYM;
    output wire BMAGYP;
    output wire BMAGZM;
    output wire BMAGZP;
    input wire BMGXM;
    input wire BMGXP;
    input wire BMGYM;
    input wire BMGYP;
    input wire BMGZM;
    input wire BMGZP;
    input wire BR1;
    input wire BR1_n;
    input wire C45R;
    input wire CA2_n;
    input wire CA4_n;
    input wire CA5_n;
    input wire CA6_n;
    input wire CAURST;
    input wire CCH11;
    input wire CCH13;
    input wire CCH14;
    output wire CCH33;
    input wire CCHG_n;
    output wire CH1109;
    output wire CH1110;
    output wire CH1111;
    output wire CH1112;
    output wire CH1305;
    output wire CH1306;
    output wire CH1308;
    output wire CH1309;
    output wire CH1401;
    output wire CH1402;
    output wire CH1403;
    output wire CH1404;
    output wire CH1405;
    output wire CH1406;
    output wire CH1407;
    output wire CH1408;
    output wire CH1409;
    output wire CH1410;
    output wire CH3310;
    output wire CH3311;
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CSG;
    input wire CXB0_n;
    input wire CXB7_n;
    output wire EMSD;
    output wire ERRST;
    input wire F04A;
    input wire F05A_n;
    input wire F05B_n;
    input wire F06B;
    input wire F07B;
    input wire F09B_n;
    input wire F10A_n;
    input wire F10B;
    output wire F5ASB0_n;
    output wire F5ASB2;
    output wire F5ASB2_n;
    output wire F5BSB2_n;
    input wire FS07A;
    input wire FS07_n;
    input wire FS10;
    input wire GATEX_n;
    input wire GATEY_n;
    input wire GATEZ_n;
    input wire GOJAM;
    input wire GTONE;
    input wire GTSET;
    input wire GTSET_n;
    output wire GYROD;
    output wire INLNKM;
    output wire INLNKP;
    input wire MOUT_n;
    output wire OTLNKM;
    input wire OVF_n;
    input wire POUT_n;
    input wire RCH11_n;
    input wire RCH13_n;
    input wire RCH14_n;
    input wire RCH33_n;
    input wire SB0_n;
    input wire SB1_n;
    input wire SB2;
    input wire SB2_n;
    input wire SHINC_n;
    input wire SIGNX;
    input wire SIGNY;
    input wire SIGNZ;
    input wire T06_n;
    output wire T1P;
    output wire T2P;
    output wire T3P;
    output wire T4P;
    output wire T5P;
    input wire T6ON_n;
    output wire T6P;
    output wire THRSTD;
    input wire UPL0;
    input wire UPL1;
    output wire UPRUPT;
    input wire WCH11_n;
    input wire WCH13_n;
    input wire WCH14_n;
    input wire WOVR_n;
    input wire XB3_n;
    input wire XB5_n;
    input wire XB6_n;
    input wire XB7_n;
    input wire XLNK0;
    input wire XLNK1;
    input wire XT3_n;
    input wire ZOUT_n;
    wire __A19_1__ALRT0;
    wire __A19_1__ALRT1;
    wire __A19_1__ALT0;
    wire __A19_1__ALT1;
    wire __A19_1__ALTSNC;
    wire __A19_1__BLKUPL;
    wire __A19_1__C45R_n;
    wire __A19_1__EMSm;
    wire __A19_1__EMSp;
    wire __A19_1__F5ASB0;
    wire __A19_1__F5BSB2;
    wire __A19_1__OTLNK0;
    wire __A19_1__OTLNK1;
    wire __A19_1__SH3MS_n;
    wire __A19_1__THRSTm;
    wire __A19_1__THRSTp;
    wire __A19_1__UPL0_n;
    wire __A19_1__UPL1_n;
    wire __A19_1__XLNK0_n;
    wire __A19_1__XLNK1_n;
    wire __A19_2__CNTRSB_n;
    wire __A19_2__F06B_n;
    wire __A19_2__F07C_n;
    wire __A19_2__F07D_n;
    wire __A19_2__F10B_n;
    wire __A19_2__F7CSB1_n;
    wire __A19_2__FF1109_n;
    wire __A19_2__FF1110_n;
    wire __A19_2__FF1111_n;
    wire __A19_2__FF1112_n;
    wire __A19_2__GYENAB;
    wire __A19_2__GYRRST;
    wire __A19_2__GYRSET;
    wire __A19_2__GYXM;
    wire __A19_2__GYXP;
    wire __A19_2__GYYM;
    wire __A19_2__GYYP;
    wire __A19_2__GYZM;
    wire __A19_2__GYZP;
    wire __A19_2__O44;
    wire __A19_2__OT1110;
    wire __A19_2__OT1111;
    wire __A19_2__OT1112;
    wire __A19_2__OUTCOM;
    wire __A19_2__RHCGO;
    wire net_U19001_Pad1;
    wire net_U19001_Pad13;
    wire net_U19001_Pad4;
    wire net_U19002_Pad11;
    wire net_U19002_Pad2;
    wire net_U19002_Pad3;
    wire net_U19002_Pad4;
    wire net_U19002_Pad5;
    wire net_U19002_Pad8;
    wire net_U19002_Pad9;
    wire net_U19003_Pad11;
    wire net_U19003_Pad6;
    wire net_U19003_Pad8;
    wire net_U19003_Pad9;
    wire net_U19004_Pad1;
    wire net_U19004_Pad10;
    wire net_U19004_Pad12;
    wire net_U19005_Pad12;
    wire net_U19006_Pad13;
    wire net_U19006_Pad3;
    wire net_U19006_Pad4;
    wire net_U19007_Pad10;
    wire net_U19007_Pad12;
    wire net_U19007_Pad6;
    wire net_U19008_Pad3;
    wire net_U19008_Pad9;
    wire net_U19009_Pad10;
    wire net_U19010_Pad1;
    wire net_U19010_Pad10;
    wire net_U19010_Pad12;
    wire net_U19010_Pad13;
    wire net_U19010_Pad4;
    wire net_U19010_Pad6;
    wire net_U19011_Pad13;
    wire net_U19011_Pad9;
    wire net_U19012_Pad1;
    wire net_U19012_Pad13;
    wire net_U19013_Pad6;
    wire net_U19014_Pad8;
    wire net_U19014_Pad9;
    wire net_U19015_Pad10;
    wire net_U19015_Pad12;
    wire net_U19015_Pad13;
    wire net_U19016_Pad10;
    wire net_U19016_Pad11;
    wire net_U19016_Pad8;
    wire net_U19016_Pad9;
    wire net_U19017_Pad10;
    wire net_U19017_Pad11;
    wire net_U19017_Pad12;
    wire net_U19017_Pad3;
    wire net_U19017_Pad9;
    wire net_U19018_Pad10;
    wire net_U19018_Pad12;
    wire net_U19018_Pad13;
    wire net_U19019_Pad1;
    wire net_U19020_Pad13;
    wire net_U19021_Pad1;
    wire net_U19021_Pad13;
    wire net_U19021_Pad3;
    wire net_U19022_Pad13;
    wire net_U19023_Pad1;
    wire net_U19024_Pad10;
    wire net_U19024_Pad8;
    wire net_U19024_Pad9;
    wire net_U19025_Pad1;
    wire net_U19025_Pad11;
    wire net_U19025_Pad4;
    wire net_U19026_Pad12;
    wire net_U19026_Pad13;
    wire net_U19027_Pad10;
    wire net_U19027_Pad4;
    wire net_U19028_Pad10;
    wire net_U19028_Pad13;
    wire net_U19029_Pad1;
    wire net_U19029_Pad10;
    wire net_U19029_Pad4;
    wire net_U19029_Pad9;
    wire net_U19030_Pad10;
    wire net_U19030_Pad11;
    wire net_U19030_Pad3;
    wire net_U19030_Pad4;
    wire net_U19030_Pad6;
    wire net_U19030_Pad8;
    wire net_U19031_Pad10;
    wire net_U19031_Pad12;
    wire net_U19031_Pad13;
    wire net_U19031_Pad4;
    wire net_U19032_Pad13;
    wire net_U19033_Pad13;
    wire net_U19034_Pad13;
    wire net_U19034_Pad3;
    wire net_U19035_Pad3;
    wire net_U19036_Pad10;
    wire net_U19036_Pad11;
    wire net_U19036_Pad12;
    wire net_U19036_Pad13;
    wire net_U19036_Pad8;
    wire net_U19037_Pad1;
    wire net_U19037_Pad10;
    wire net_U19038_Pad1;
    wire net_U19038_Pad10;
    wire net_U19039_Pad1;
    wire net_U19039_Pad13;
    wire net_U19040_Pad1;
    wire net_U19040_Pad13;
    wire net_U19040_Pad3;
    wire net_U19041_Pad1;
    wire net_U19041_Pad13;
    wire net_U19042_Pad13;
    wire net_U19042_Pad3;
    wire net_U19043_Pad1;
    wire net_U19043_Pad3;
    wire net_U19044_Pad10;
    wire net_U19044_Pad11;
    wire net_U19044_Pad8;
    wire net_U19044_Pad9;
    wire net_U19046_Pad13;
    wire net_U19047_Pad11;
    wire net_U19047_Pad13;
    wire net_U19047_Pad2;
    wire net_U19047_Pad3;
    wire net_U19047_Pad9;
    wire net_U19049_Pad10;
    wire net_U19049_Pad13;
    wire net_U19050_Pad10;
    wire net_U19050_Pad12;
    wire net_U19050_Pad13;
    wire net_U19051_Pad1;
    wire net_U19051_Pad10;
    wire net_U19051_Pad2;
    wire net_U19051_Pad3;
    wire net_U19052_Pad10;
    wire net_U19052_Pad13;
    wire net_U19053_Pad8;
    wire net_U19053_Pad9;
    wire net_U19055_Pad6;
    wire net_U19055_Pad8;
    wire net_U19056_Pad10;
    wire net_U19056_Pad12;
    wire net_U19056_Pad13;
    wire net_U19056_Pad4;
    wire net_U19057_Pad10;
    wire net_U19057_Pad12;
    wire net_U19057_Pad13;
    wire net_U19057_Pad4;
    wire net_U19057_Pad6;
    wire net_U19057_Pad9;
    wire net_U19059_Pad12;
    wire net_U19059_Pad6;
    wire net_U19059_Pad8;
    wire net_U19060_Pad1;
    wire net_U19060_Pad10;
    wire net_U19060_Pad4;

    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19001(net_U19001_Pad1, CA6_n, CXB0_n, net_U19001_Pad4, SHINC_n, T06_n, GND, net_U19001_Pad4, net_U19001_Pad13, __A19_1__SH3MS_n, __A19_1__SH3MS_n, CSG, net_U19001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U19002(net_U19001_Pad1, net_U19002_Pad2, net_U19002_Pad3, net_U19002_Pad4, net_U19002_Pad5, __A19_1__ALTSNC, GND, net_U19002_Pad8, net_U19002_Pad9, __A19_1__OTLNK0, net_U19002_Pad11, F5ASB0_n, __A19_1__F5ASB0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19003(BR1, __A19_1__SH3MS_n, net_U19002_Pad2, __A19_1__SH3MS_n, BR1_n, net_U19003_Pad6, GND, net_U19003_Pad8, net_U19003_Pad9, CCH14, net_U19003_Pad11, net_U19002_Pad3, net_U19002_Pad2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19004(net_U19004_Pad1, CHWL02_n, WCH14_n, net_U19004_Pad12, net_U19004_Pad1, net_U19004_Pad10, GND, net_U19004_Pad12, CCH14, net_U19004_Pad10, RCH14_n, net_U19004_Pad12, CH1402, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19005(__A19_1__ALT0, net_U19002_Pad4, net_U19004_Pad10, __A19_1__ALT1, net_U19004_Pad10, net_U19005_Pad12, GND, net_U19002_Pad4, net_U19004_Pad12, __A19_1__ALRT0, net_U19004_Pad12, net_U19005_Pad12, __A19_1__ALRT1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19006(net_U19005_Pad12, net_U19003_Pad6, net_U19006_Pad3, net_U19006_Pad4, WCH14_n, CHWL03_n, GND, net_U19006_Pad4, net_U19003_Pad8, net_U19003_Pad9, net_U19003_Pad8, net_U19003_Pad11, net_U19006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19007(CH1403, RCH14_n, net_U19006_Pad13, net_U19007_Pad12, net_U19007_Pad10, net_U19007_Pad6, GND, net_U19003_Pad9, GTSET_n, net_U19007_Pad10, F5ASB2_n, net_U19007_Pad12, net_U19006_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19008(net_U19007_Pad12, GOJAM, net_U19008_Pad3, GTSET, GOJAM, net_U19003_Pad11, GND, net_U19002_Pad5, net_U19008_Pad9, net_U19003_Pad11, net_U19007_Pad6, net_U19007_Pad6, GTONE, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U19009(net_U19008_Pad3, net_U19006_Pad3, net_U19003_Pad11, ALTM, F5ASB0_n, net_U19008_Pad3, GND, net_U19003_Pad11, net_U19008_Pad9, net_U19009_Pad10, net_U19009_Pad10, GTONE, net_U19008_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19010(net_U19010_Pad1, CHWL01_n, WCH14_n, net_U19010_Pad4, net_U19010_Pad1, net_U19010_Pad6, GND, GTSET_n, net_U19010_Pad4, net_U19010_Pad10, net_U19010_Pad10, net_U19010_Pad12, net_U19010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19011(net_U19010_Pad4, CCH14, net_U19010_Pad13, GTONE, GOJAM, net_U19010_Pad12, GND, net_U19011_Pad13, net_U19011_Pad9, GTSET, GOJAM, net_U19010_Pad6, net_U19011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19012(net_U19012_Pad1, F5ASB2_n, net_U19010_Pad13, net_U19011_Pad9, net_U19012_Pad1, net_U19011_Pad13, GND, F5ASB0_n, net_U19011_Pad9, OTLNKM, net_U19010_Pad6, net_U19011_Pad13, net_U19012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19013(CH1401, net_U19012_Pad13, RCH14_n, net_U19002_Pad11, net_U19012_Pad1, net_U19013_Pad6, GND, CA5_n, CXB7_n, net_U19002_Pad9, SB0_n, F05A_n, __A19_1__F5ASB0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19014(BR1_n, __A19_1__SH3MS_n, net_U19002_Pad8, __A19_1__SH3MS_n, BR1, __A19_1__OTLNK1, GND, net_U19014_Pad8, net_U19014_Pad9, __A19_1__UPL0_n, __A19_1__BLKUPL, net_U19013_Pad6, net_U19002_Pad8, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19015(F5ASB2, F05A_n, SB2_n, __A19_1__F5BSB2, SB2_n, F05B_n, GND, __A19_1__XLNK0_n, net_U19015_Pad12, net_U19015_Pad10, __A19_1__XLNK1_n, net_U19015_Pad12, net_U19015_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U19016(F5ASB2, F5ASB2_n, __A19_1__F5BSB2, F5BSB2_n, C45R, __A19_1__C45R_n, GND, net_U19016_Pad8, net_U19016_Pad9, net_U19016_Pad10, net_U19016_Pad11, __A19_1__UPL0_n, UPL0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19017(__A19_1__BLKUPL, net_U19014_Pad9, net_U19017_Pad3, net_U19017_Pad10, net_U19017_Pad11, INLNKM, GND, INLNKP, net_U19017_Pad9, net_U19017_Pad10, net_U19017_Pad11, net_U19017_Pad12, __A19_1__UPL1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U19018(net_U19017_Pad3, net_U19014_Pad8, net_U19015_Pad10, net_U19017_Pad9, net_U19017_Pad12, net_U19015_Pad13, GND, __A19_1__C45R_n, net_U19018_Pad13, net_U19018_Pad10, net_U19018_Pad10, net_U19018_Pad12, net_U19018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U19019(net_U19019_Pad1, net_U19014_Pad8, net_U19017_Pad12, net_U19015_Pad10, net_U19015_Pad13,  , GND,  , CA2_n, XB5_n, WOVR_n, OVF_n, T2P, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19020(net_U19018_Pad12, net_U19018_Pad10, net_U19017_Pad11, net_U19017_Pad11, net_U19018_Pad12, F04A, GND, BR1_n, __A19_1__C45R_n, UPRUPT, net_U19018_Pad12, net_U19019_Pad1, net_U19020_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19021(net_U19021_Pad1, net_U19020_Pad13, net_U19021_Pad3, CH3311, net_U19021_Pad3, RCH33_n, GND, RCH33_n, __A19_1__BLKUPL, CH3310, CHWL05_n, WCH13_n, net_U19021_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19022(net_U19015_Pad12, net_U19021_Pad13, net_U19014_Pad9, net_U19014_Pad9, net_U19015_Pad12, CCH13, GND, net_U19015_Pad12, RCH13_n, CH1305, WCH13_n, CHWL06_n, net_U19022_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19023(net_U19023_Pad1, net_U19022_Pad13, net_U19017_Pad10, net_U19017_Pad10, net_U19023_Pad1, CCH13, GND, net_U19023_Pad1, RCH13_n, CH1306, CA5_n, XB5_n, net_U19016_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19024(net_U19021_Pad1, CCH33, CCHG_n, XT3_n, XB3_n, CCH33, GND, net_U19024_Pad8, net_U19024_Pad9, net_U19024_Pad10, CCH14, net_U19021_Pad3, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19025(net_U19025_Pad1, net_U19016_Pad8, POUT_n, net_U19025_Pad4, net_U19016_Pad8, MOUT_n, GND, net_U19016_Pad8, ZOUT_n, net_U19024_Pad10, net_U19025_Pad11, net_U19024_Pad8, net_U19024_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19026(net_U19025_Pad11, WCH14_n, CHWL04_n, CH1404, RCH14_n, net_U19024_Pad9, GND, net_U19024_Pad9, F5ASB2_n, THRSTD, net_U19025_Pad1, net_U19026_Pad12, net_U19026_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19027(net_U19026_Pad12, net_U19026_Pad13, net_U19024_Pad9, net_U19027_Pad4, net_U19025_Pad4, net_U19027_Pad10, GND, net_U19027_Pad4, net_U19024_Pad9, net_U19027_Pad10, net_U19026_Pad13, F5ASB0_n, __A19_1__THRSTp, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19028(__A19_1__THRSTm, net_U19027_Pad4, F5ASB0_n, net_U19016_Pad11, CA5_n, XB6_n, GND, net_U19016_Pad10, POUT_n, net_U19028_Pad10, WCH14_n, CHWL05_n, net_U19028_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19029(net_U19029_Pad1, net_U19016_Pad10, MOUT_n, net_U19029_Pad4, net_U19016_Pad10, ZOUT_n, GND, net_U19028_Pad13, net_U19029_Pad9, net_U19029_Pad10, RCH14_n, net_U19029_Pad10, CH1405, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19030(net_U19029_Pad10, net_U19029_Pad4, net_U19030_Pad3, net_U19030_Pad4, CCH14, net_U19030_Pad6, GND, net_U19030_Pad8, SB1_n, net_U19030_Pad10, net_U19030_Pad11, net_U19029_Pad9, CCH14, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19031(EMSD, net_U19029_Pad10, F5ASB2_n, net_U19031_Pad4, net_U19028_Pad10, net_U19031_Pad10, GND, net_U19031_Pad4, net_U19029_Pad10, net_U19031_Pad10, net_U19029_Pad1, net_U19031_Pad12, net_U19031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19032(net_U19031_Pad12, net_U19031_Pad13, net_U19029_Pad10, __A19_1__EMSp, net_U19031_Pad4, F5ASB0_n, GND, net_U19031_Pad13, F5ASB0_n, __A19_1__EMSm, CHWL09_n, WCH11_n, net_U19032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U19033(BLKUPL_n, __A19_1__BLKUPL, UPL1, __A19_1__UPL1_n, XLNK0, __A19_1__XLNK0_n, GND, __A19_1__XLNK1_n, XLNK1, __A19_2__OUTCOM, __A19_2__FF1109_n, ERRST, net_U19033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19034(__A19_2__FF1109_n, net_U19032_Pad13, net_U19034_Pad3, net_U19034_Pad3, __A19_2__FF1109_n, CCH11, GND, RCH11_n, __A19_2__FF1109_n, CH1109, CHWL10_n, WCH11_n, net_U19034_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19035(__A19_2__FF1110_n, net_U19034_Pad13, net_U19035_Pad3, net_U19035_Pad3, __A19_2__FF1110_n, CCH11, GND, CAURST, net_U19034_Pad13, net_U19033_Pad13, RCH11_n, __A19_2__FF1110_n, CH1110, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U19036(__A19_2__FF1110_n, __A19_2__OT1110, __A19_2__FF1111_n, __A19_2__OT1111, __A19_2__FF1112_n, __A19_2__OT1112, GND, net_U19036_Pad8, net_U19030_Pad8, net_U19036_Pad10, net_U19036_Pad11, net_U19036_Pad12, net_U19036_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19037(net_U19037_Pad1, CHWL11_n, WCH11_n, __A19_2__FF1111_n, net_U19037_Pad1, net_U19037_Pad10, GND, __A19_2__FF1111_n, CCH11, net_U19037_Pad10, RCH11_n, __A19_2__FF1111_n, CH1111, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19038(net_U19038_Pad1, CHWL12_n, WCH11_n, __A19_2__FF1112_n, net_U19038_Pad1, net_U19038_Pad10, GND, __A19_2__FF1112_n, CCH11, net_U19038_Pad10, RCH11_n, __A19_2__FF1112_n, CH1112, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19039(net_U19039_Pad1, CHWL10_n, WCH14_n, net_U19030_Pad3, net_U19039_Pad1, net_U19030_Pad6, GND, RCH14_n, net_U19030_Pad3, CH1410, CHWL09_n, WCH14_n, net_U19039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19040(net_U19040_Pad1, net_U19039_Pad13, net_U19040_Pad3, net_U19040_Pad3, net_U19040_Pad1, CCH14, GND, RCH14_n, net_U19040_Pad1, CH1409, CHWL08_n, WCH14_n, net_U19040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19041(net_U19041_Pad1, net_U19040_Pad13, net_U19030_Pad10, net_U19030_Pad10, net_U19041_Pad1, CCH14, GND, RCH14_n, net_U19041_Pad1, CH1408, CHWL07_n, WCH14_n, net_U19041_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19042(net_U19030_Pad11, net_U19041_Pad13, net_U19042_Pad3, net_U19042_Pad3, net_U19030_Pad11, CCH14, GND, RCH14_n, net_U19030_Pad11, CH1407, CHWL06_n, WCH14_n, net_U19042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19043(net_U19043_Pad1, net_U19042_Pad13, net_U19043_Pad3, net_U19043_Pad3, net_U19043_Pad1, CCH14, GND, RCH14_n, net_U19043_Pad1, CH1406, net_U19030_Pad3, F5ASB2_n, GYROD, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19044(SB1_n, net_U19042_Pad3, SB1_n, net_U19041_Pad1, net_U19030_Pad11, net_U19036_Pad13, GND, net_U19044_Pad8, net_U19044_Pad9, net_U19044_Pad10, net_U19044_Pad11, net_U19036_Pad11, net_U19041_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19045(__A19_2__GYENAB, SB1_n, net_U19043_Pad1, __A19_2__GYXP, net_U19040_Pad3, net_U19036_Pad8, GND, net_U19036_Pad8, net_U19040_Pad1, __A19_2__GYXM, net_U19040_Pad3, net_U19036_Pad10, __A19_2__GYYP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19046(__A19_2__GYYM, net_U19036_Pad10, net_U19040_Pad1, __A19_2__GYZP, net_U19040_Pad3, net_U19036_Pad12, GND, net_U19036_Pad12, net_U19040_Pad1, __A19_2__GYZM, CA4_n, XB7_n, net_U19046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0) U19047(net_U19046_Pad13, net_U19047_Pad2, net_U19047_Pad3, __A19_2__O44, F06B, __A19_2__F06B_n, GND, __A19_2__F07D_n, net_U19047_Pad9, __A19_2__F07C_n, net_U19047_Pad11, __A19_2__F7CSB1_n, net_U19047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19048(net_U19044_Pad10, POUT_n, net_U19047_Pad2, net_U19044_Pad11, MOUT_n, net_U19047_Pad2, GND, ZOUT_n, net_U19047_Pad2, net_U19030_Pad4, net_U19030_Pad3, net_U19044_Pad8, net_U19044_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19049(__A19_2__GYRRST, F5ASB2_n, net_U19044_Pad9, __A19_2__GYRSET, F5ASB2_n, net_U19044_Pad8, GND, CHWL08_n, WCH13_n, net_U19049_Pad10, net_U19049_Pad10, net_U19047_Pad3, net_U19049_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19050(net_U19047_Pad3, net_U19049_Pad13, CCH13, CH1308, RCH13_n, net_U19049_Pad13, GND, WCH13_n, CHWL09_n, net_U19050_Pad10, net_U19050_Pad10, net_U19050_Pad12, net_U19050_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19051(net_U19051_Pad1, net_U19051_Pad2, net_U19051_Pad3, CH1309, RCH13_n, net_U19050_Pad13, GND, net_U19050_Pad13, __A19_2__F07D_n, net_U19051_Pad10, FS07_n, __A19_2__F06B_n, net_U19047_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19052(net_U19047_Pad11, __A19_2__F06B_n, FS07A, net_U19047_Pad13, __A19_2__F07C_n, SB1_n, GND, net_U19051_Pad10, net_U19052_Pad13, net_U19052_Pad10, net_U19052_Pad10, F07B, net_U19052_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19053(SB2_n, net_U19052_Pad10, net_U19050_Pad13, CCH13, __A19_2__RHCGO, net_U19050_Pad12, GND, net_U19053_Pad8, net_U19053_Pad9, __A19_2__F07C_n, SB0_n, __A19_2__RHCGO, __A19_2__F07C_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U19054(net_U19052_Pad13, net_U19053_Pad9, SB2, __A19_2__CNTRSB_n, F10B, __A19_2__F10B_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19055(SIGNX, net_U19053_Pad9, SIGNY, net_U19053_Pad9, __A19_2__F7CSB1_n, net_U19055_Pad6, GND, net_U19055_Pad8, SIGNZ, net_U19053_Pad9, __A19_2__F7CSB1_n, net_U19051_Pad2, __A19_2__F7CSB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19056(net_U19051_Pad3, net_U19051_Pad1, net_U19053_Pad8, net_U19056_Pad4, net_U19055_Pad6, net_U19056_Pad10, GND, net_U19056_Pad4, net_U19053_Pad8, net_U19056_Pad10, net_U19055_Pad8, net_U19056_Pad12, net_U19056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19057(net_U19056_Pad12, net_U19056_Pad13, net_U19053_Pad8, net_U19057_Pad4, BMGXP, net_U19057_Pad6, GND, BMGXM, net_U19057_Pad9, net_U19057_Pad10, BMGYP, net_U19057_Pad12, net_U19057_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19058(F5ASB2_n, net_U19051_Pad1, F5ASB2_n, net_U19051_Pad3, GATEX_n, net_U19057_Pad9, GND, net_U19057_Pad12, F5ASB2_n, net_U19056_Pad4, GATEY_n, net_U19057_Pad6, GATEX_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19059(F5ASB2_n, net_U19056_Pad10, F5ASB2_n, net_U19056_Pad13, GATEZ_n, net_U19059_Pad6, GND, net_U19059_Pad8, F5ASB2_n, net_U19056_Pad12, GATEZ_n, net_U19059_Pad12, GATEY_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19060(net_U19060_Pad1, BMGYM, net_U19059_Pad12, net_U19060_Pad4, BMGZP, net_U19059_Pad6, GND, BMGZM, net_U19059_Pad8, net_U19060_Pad10, __A19_2__O44, net_U19057_Pad4, BMAGXP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19061(BMAGXM, __A19_2__O44, net_U19057_Pad10, BMAGYP, __A19_2__O44, net_U19057_Pad13, GND, __A19_2__O44, net_U19060_Pad1, BMAGYM, __A19_2__O44, net_U19060_Pad4, BMAGZP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19062(BMAGZM, __A19_2__O44, net_U19060_Pad10, T1P, __A19_2__CNTRSB_n, __A19_2__F10B_n, GND, __A19_2__F10B_n, __A19_2__CNTRSB_n, T3P, F10A_n, __A19_2__CNTRSB_n, T5P, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19063(FS10, F09B_n, __A19_2__F06B_n, T6ON_n, __A19_2__CNTRSB_n, T6P, GND,  ,  ,  ,  , T4P, __A19_2__CNTRSB_n, p4VSW, SIM_RST, SIM_CLK);
endmodule