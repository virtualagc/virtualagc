// Verilog testbench created by dumbTestbench.py
`timescale 100ns / 1ns

module agc;

`include "2005250-/tb.v"

reg ALTM = 0, BMAGXM = 0, BMAGXP = 0, BMAGYM = 0, BMAGYP = 0, BMAGZM = 0,
  BMAGZP = 0, C24A = 0, C25A = 0, C26A = 0, C27A = 0, C30A = 0, C31A = 0,
  C32A = 0, C33A = 0, C34A = 0, C35A = 0, C36A = 0, C37A = 0, C40A = 0,
  C41A = 0, C50A = 0, C51A = 0, C52A = 0, C53A = 0, C54A = 0, C55A = 0,
  CA6_ = 0, CG13 = 0, CG23 = 0, CGA21 = 0, CT = 0, CXB2_ = 0, CXB3_ = 0,
  CXB4_ = 0, CXB7_ = 0, DOSCAL = 0, EMSD = 0, FS17 = 0, GNHNC = 0, GOJAM = 0,
  GYROD = 0, INLNKM = 0, INLNKP = 0, MLDCH = 0, MLOAD = 0, MNHNC = 0, MRDCH = 0,
  MREAD = 0, NISQL_ = 0, OCTAD4 = 0, OCTAD5 = 0, OTLNKM = 0, PHS2_ = 0,
  PHS3_ = 0, PHS4_ = 0, PSEUDO = 0, RNRADM = 0, RNRADP = 0, RQ = 0, RSCT_ = 0,
  ST0_ = 0, ST1_ = 0, STD2 = 0, T02_ = 0, T07_ = 0, T10_ = 0, T11_ = 0,
  T12A = 0, T12_ = 0, XB0 = 0, XB5 = 0, XB6 = 0;

wire BKTF_, C42A, C42M, C42P, C42R, C43A, C43M, C43P, C43R, C44A, C44M,
  C44P, C44R, C45A, C45M, C45P, C45R, C46A, C46M, C46P, C46R, C47A, C47R,
  C56A, C56R, C57A, C57R, C60A, C60R, CA4_, CA5_, CAD1, CAD2, CAD3, CAD4,
  CAD5, CAD6, CG15, CG16, CG26, CHINC, CHINC_, CTROR, CTROR_, CXB0_, CXB5_,
  CXB6_, DINC, DINCNC_, DINC_, FETCH0, FETCH0_, FETCH1, INCSET_, INKBT1,
  INKL, INKL_, INOTLD, INOTRD, MINKL, MON_, MONpCH, MREQIN, RQ_, RSSB,
  SCAS17, SHANC, SHANC_, SHINC, SHINC_, STFET1_, STORE1, STORE1_, d30SUM,
  d32004K, d50SUM;

A21 iA21 (
  rst, ALTM, BMAGXM, BMAGXP, BMAGYM, BMAGYP, BMAGZM, BMAGZP, C24A, C25A,
  C26A, C27A, C30A, C31A, C32A, C33A, C34A, C35A, C36A, C37A, C40A, C41A,
  C50A, C51A, C52A, C53A, C54A, C55A, CA6_, CG13, CG23, CGA21, CT, CXB2_,
  CXB3_, CXB4_, CXB7_, DOSCAL, EMSD, FS17, GNHNC, GOJAM, GYROD, INLNKM, INLNKP,
  MLDCH, MLOAD, MNHNC, MRDCH, MREAD, NISQL_, OCTAD4, OCTAD5, OTLNKM, PHS2_,
  PHS3_, PHS4_, PSEUDO, RNRADM, RNRADP, RQ, RSCT_, ST0_, ST1_, STD2, T02_,
  T07_, T10_, T11_, T12A, T12_, XB0, XB5, XB6, BKTF_, C42A, C43A, C44A, C45A,
  C45M, C45P, C46A, C46M, C46P, C47A, C56A, C57A, C60A, CA4_, CA5_, CG15,
  CG16, CHINC, CHINC_, CTROR_, CXB0_, CXB5_, CXB6_, DINC, INCSET_, INKBT1,
  INOTLD, INOTRD, MINKL, MREQIN, RSSB, SCAS17, d32004K, C42M, C42P, C42R,
  C43M, C43P, C43R, C44M, C44P, C44R, C45R, C46R, C47R, C56R, C57R, C60R,
  CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CG26, CTROR, DINCNC_, DINC_, FETCH0,
  FETCH0_, FETCH1, INKL, INKL_, MON_, MONpCH, RQ_, SHANC, SHANC_, SHINC,
  SHINC_, STFET1_, STORE1, STORE1_, d30SUM, d50SUM
);

endmodule
