`timescale 1ns/1ps
`default_nettype none

module rupt_service(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, T10, S10, S10_n, S11_n, S12_n, WL01_n, WL02_n, WL03_n, WL09_n, WL10_n, WL11_n, WL12_n, WL13_n, WL14_n, WL16_n, SUMA01_n, SUMB01_n, SUMA02_n, SUMB02_n, SUMA03_n, SUMB03_n, SUMA11_n, SUMB11_n, SUMA12_n, SUMB12_n, SUMA13_n, SUMB13_n, SUMA14_n, SUMB14_n, SUMA16_n, SUMB16_n, XB0_n, XB1_n, XB4_n, XB6_n, XB7_n, XT0_n, XT1_n, XT2_n, XT3_n, XT4_n, XT5_n, E5, E6, E7_n, STRGAT, CEBG, CFBG, OVF_n, R6, RB1F, RBBEG_n, REBG_n, RFBG_n, RRPA, RSTRT, U2BBKG_n, WBBEG_n, WEBG_n, WFBG_n, WOVR_n, ZOUT_n, DLKPLS, HNDRPT, KRPT, KYRPT1, KYRPT2, RADRPT, UPRUPT, CA2_n, CA3_n, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, MKRPT, EB9, EB10, EB11_n, RL01_n, RL02_n, RL03_n, RL04_n, RL05_n, RL06_n, RL09_n, RL10_n, RL11_n, RL12_n, RL13_n, RL14_n, RL15_n, RL16_n, RUPTOR_n, ROPER, ROPES, ROPET, HIMOD, LOMOD, STR19, STR210, STR311, STR412, STR14, STR58, STR912, T6RPT, DRPRST, STRT2);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire CA2_n;
    input wire CA3_n;
    input wire CAD1;
    input wire CAD2;
    input wire CAD3;
    input wire CAD4;
    input wire CAD5;
    input wire CAD6;
    input wire CEBG;
    input wire CFBG;
    input wire DLKPLS;
    output wire DRPRST;
    input wire E5;
    input wire E6;
    input wire E7_n;
    output wire EB10;
    output wire EB11_n;
    output wire EB9;
    input wire GOJAM;
    output wire HIMOD;
    input wire HNDRPT;
    input wire KRPT;
    input wire KYRPT1;
    input wire KYRPT2;
    output wire LOMOD;
    input wire MKRPT;
    input wire OVF_n;
    input wire R6;
    input wire RADRPT;
    input wire RB1F;
    input wire RBBEG_n;
    input wire REBG_n;
    input wire RFBG_n;
    output wire RL01_n; //FPGA#wand
    output wire RL02_n; //FPGA#wand
    output wire RL03_n; //FPGA#wand
    output wire RL04_n; //FPGA#wand
    output wire RL05_n; //FPGA#wand
    output wire RL06_n; //FPGA#wand
    output wire RL09_n; //FPGA#wand
    output wire RL10_n; //FPGA#wand
    output wire RL11_n; //FPGA#wand
    output wire RL12_n; //FPGA#wand
    output wire RL13_n; //FPGA#wand
    output wire RL14_n; //FPGA#wand
    output wire RL15_n; //FPGA#wand
    output wire RL16_n; //FPGA#wand
    output wire ROPER;
    output wire ROPES;
    output wire ROPET;
    input wire RRPA;
    input wire RSTRT;
    output wire RUPTOR_n;
    input wire S10;
    input wire S10_n;
    input wire S11_n;
    input wire S12_n;
    output wire STR14;
    output wire STR19;
    output wire STR210;
    output wire STR311;
    output wire STR412;
    output wire STR58;
    output wire STR912;
    input wire STRGAT;
    input wire STRT2;
    input wire SUMA01_n;
    input wire SUMA02_n;
    input wire SUMA03_n;
    input wire SUMA11_n;
    input wire SUMA12_n;
    input wire SUMA13_n;
    input wire SUMA14_n;
    input wire SUMA16_n;
    input wire SUMB01_n;
    input wire SUMB02_n;
    input wire SUMB03_n;
    input wire SUMB11_n;
    input wire SUMB12_n;
    input wire SUMB13_n;
    input wire SUMB14_n;
    input wire SUMB16_n;
    input wire T10;
    output wire T6RPT;
    input wire U2BBKG_n;
    input wire UPRUPT;
    input wire WBBEG_n;
    input wire WEBG_n;
    input wire WFBG_n;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL16_n;
    input wire WOVR_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB4_n;
    input wire XB6_n;
    input wire XB7_n;
    input wire XT0_n;
    input wire XT1_n;
    input wire XT2_n;
    input wire XT3_n;
    input wire XT4_n;
    input wire XT5_n;
    input wire ZOUT_n;
    wire __A15_1__BBK1;
    wire __A15_1__BBK2;
    wire __A15_1__BBK3;
    wire __A15_1__BK16;
    wire __A15_1__DNRPTA;
    wire __A15_1__EB10_n;
    wire __A15_1__EB11;
    wire __A15_1__EB9_n;
    wire __A15_1__F11;
    wire __A15_1__F11_n;
    wire __A15_1__F12;
    wire __A15_1__F12_n;
    wire __A15_1__F13;
    wire __A15_1__F13_n;
    wire __A15_1__F14;
    wire __A15_1__F14_n;
    wire __A15_1__F15;
    wire __A15_1__F15_n;
    wire __A15_1__F16;
    wire __A15_1__F16_n;
    wire __A15_1__FB11;
    wire __A15_1__FB11_n;
    wire __A15_1__FB12;
    wire __A15_1__FB12_n;
    wire __A15_1__FB13;
    wire __A15_1__FB13_n;
    wire __A15_1__FB14;
    wire __A15_1__FB14_n;
    wire __A15_1__FB16;
    wire __A15_1__FB16_n;
    wire __A15_1__KRPTA_n;
    wire __A15_1__PRPOR1;
    wire __A15_1__PRPOR2;
    wire __A15_1__PRPOR3;
    wire __A15_1__PRPOR4;
    wire __A15_1__RPTA12;
    wire __A15_1__RPTAD6;
    wire __A15_1__RRPA1_n;
    wire __A15_2__036H;
    wire __A15_2__036L;
    wire __A15_2__147H;
    wire __A15_2__147L;
    wire __A15_2__2510H;
    wire __A15_2__2510L;
    wire __A15_2__KY1RST;
    wire __A15_2__KY2RST;
    wire __A15_2__NE00;
    wire __A15_2__NE01;
    wire __A15_2__NE012_n;
    wire __A15_2__NE02;
    wire __A15_2__NE03;
    wire __A15_2__NE036_n;
    wire __A15_2__NE04;
    wire __A15_2__NE05;
    wire __A15_2__NE06;
    wire __A15_2__NE07;
    wire __A15_2__NE10;
    wire __A15_2__NE147_n;
    wire __A15_2__NE2510_n;
    wire __A15_2__NE345_n;
    wire __A15_2__NE6710_n;
    wire __A15_2__RPTAD3;
    wire __A15_2__RPTAD4;
    wire __A15_2__RPTAD5;
    wire net_R15001_Pad2; //FPGA#wand
    wire net_R15002_Pad2; //FPGA#wand
    wire net_U15001_Pad1;
    wire net_U15001_Pad13;
    wire net_U15002_Pad2;
    wire net_U15002_Pad8;
    wire net_U15003_Pad10;
    wire net_U15003_Pad11;
    wire net_U15003_Pad12;
    wire net_U15003_Pad13;
    wire net_U15003_Pad2;
    wire net_U15003_Pad4;
    wire net_U15003_Pad5;
    wire net_U15003_Pad6;
    wire net_U15003_Pad8;
    wire net_U15003_Pad9;
    wire net_U15004_Pad11;
    wire net_U15004_Pad13;
    wire net_U15005_Pad10;
    wire net_U15005_Pad9;
    wire net_U15007_Pad13;
    wire net_U15007_Pad4;
    wire net_U15008_Pad12;
    wire net_U15009_Pad1;
    wire net_U15009_Pad10;
    wire net_U15009_Pad12;
    wire net_U15010_Pad12;
    wire net_U15010_Pad8;
    wire net_U15011_Pad1;
    wire net_U15011_Pad4;
    wire net_U15012_Pad10;
    wire net_U15012_Pad11;
    wire net_U15012_Pad9;
    wire net_U15014_Pad10;
    wire net_U15014_Pad6;
    wire net_U15014_Pad9;
    wire net_U15015_Pad10;
    wire net_U15015_Pad13;
    wire net_U15016_Pad11;
    wire net_U15016_Pad13;
    wire net_U15016_Pad5;
    wire net_U15016_Pad9;
    wire net_U15018_Pad13;
    wire net_U15020_Pad3;
    wire net_U15021_Pad4;
    wire net_U15022_Pad10;
    wire net_U15022_Pad11;
    wire net_U15022_Pad13;
    wire net_U15022_Pad3;
    wire net_U15022_Pad4;
    wire net_U15022_Pad8;
    wire net_U15022_Pad9;
    wire net_U15023_Pad10;
    wire net_U15023_Pad6;
    wire net_U15023_Pad8;
    wire net_U15023_Pad9;
    wire net_U15024_Pad12;
    wire net_U15024_Pad4;
    wire net_U15024_Pad6;
    wire net_U15024_Pad8;
    wire net_U15027_Pad4;
    wire net_U15028_Pad3;
    wire net_U15028_Pad5;
    wire net_U15028_Pad6;
    wire net_U15029_Pad10;
    wire net_U15029_Pad11;
    wire net_U15029_Pad12;
    wire net_U15029_Pad13;
    wire net_U15029_Pad4;
    wire net_U15029_Pad5;
    wire net_U15029_Pad6;
    wire net_U15029_Pad8;
    wire net_U15029_Pad9;
    wire net_U15030_Pad5;
    wire net_U15031_Pad5;
    wire net_U15032_Pad5;
    wire net_U15033_Pad1;
    wire net_U15033_Pad10;
    wire net_U15033_Pad13;
    wire net_U15033_Pad3;
    wire net_U15033_Pad4;
    wire net_U15033_Pad6;
    wire net_U15034_Pad11;
    wire net_U15034_Pad8;
    wire net_U15035_Pad11;
    wire net_U15037_Pad10;
    wire net_U15037_Pad13;
    wire net_U15037_Pad3;
    wire net_U15038_Pad1;
    wire net_U15038_Pad10;
    wire net_U15038_Pad8;
    wire net_U15039_Pad11;
    wire net_U15039_Pad13;
    wire net_U15039_Pad3;
    wire net_U15039_Pad5;
    wire net_U15039_Pad9;
    wire net_U15041_Pad1;
    wire net_U15044_Pad10;
    wire net_U15044_Pad12;
    wire net_U15044_Pad4;
    wire net_U15044_Pad6;
    wire net_U15044_Pad8;
    wire net_U15048_Pad1;
    wire net_U15048_Pad10;
    wire net_U15048_Pad4;
    wire net_U15049_Pad10;
    wire net_U15049_Pad12;
    wire net_U15049_Pad2;
    wire net_U15049_Pad4;
    wire net_U15049_Pad6;
    wire net_U15049_Pad8;
    wire net_U15052_Pad9;
    wire net_U15053_Pad11;
    wire net_U15053_Pad3;
    wire net_U15053_Pad9;
    wire net_U15057_Pad13;
    wire net_U15058_Pad6;

    pullup R15001(net_R15001_Pad2);
    pullup R15002(net_R15002_Pad2);
    U74HC02 U15001(net_U15001_Pad1, WL16_n, WFBG_n, __A15_1__FB16, __A15_1__FB16_n, CFBG, GND, __A15_1__FB16_n, RFBG_n, __A15_1__BK16, WL14_n, WFBG_n, net_U15001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U15002(net_U15001_Pad1, net_U15002_Pad2, SUMA16_n, U2BBKG_n, SUMB16_n, net_U15002_Pad2, GND, net_U15002_Pad8, SUMA14_n, U2BBKG_n, SUMB14_n, __A15_1__FB16_n, __A15_1__FB16, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15003(__A15_1__BK16, net_U15003_Pad2, __A15_1__BK16, net_U15003_Pad4, net_U15003_Pad5, net_U15003_Pad6, GND, net_U15003_Pad8, net_U15003_Pad9, net_U15003_Pad10, net_U15003_Pad11, net_U15003_Pad12, net_U15003_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15004(net_U15003_Pad2, RL16_n, net_U15003_Pad4, RL15_n, net_U15003_Pad6, RL14_n, GND, RL13_n, net_U15003_Pad8, RL12_n, net_U15004_Pad11, RL11_n, net_U15004_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1) U15005(net_U15001_Pad13, net_U15002_Pad8, SUMA13_n, U2BBKG_n, SUMB13_n, net_U15005_Pad10, GND, __A15_1__FB13_n, net_U15005_Pad9, net_U15005_Pad10, __A15_1__FB13, __A15_1__FB14_n, __A15_1__FB14, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15006(__A15_1__FB14, __A15_1__FB14_n, CFBG, net_U15003_Pad5, __A15_1__FB14_n, RFBG_n, GND, WL13_n, WFBG_n, net_U15005_Pad9, __A15_1__FB13_n, CFBG, __A15_1__FB13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15007(net_U15003_Pad9, __A15_1__FB13_n, RFBG_n, net_U15007_Pad4, WL12_n, WFBG_n, GND, __A15_1__FB12_n, CFBG, __A15_1__FB12, __A15_1__FB12_n, RFBG_n, net_U15007_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U15008(SUMA12_n, U2BBKG_n, net_U15007_Pad4, net_U15008_Pad12, __A15_1__FB12, __A15_1__FB12_n, GND, net_U15004_Pad11, RSTRT, net_U15007_Pad13, __A15_1__RPTA12, net_U15008_Pad12, SUMB12_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15009(net_U15009_Pad1, WFBG_n, WL11_n, __A15_1__FB11, __A15_1__FB11_n, CFBG, GND, __A15_1__FB11_n, RFBG_n, net_U15009_Pad10, net_U15009_Pad10, net_U15009_Pad12, net_U15004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U15010(SUMA11_n, U2BBKG_n, net_U15009_Pad1, net_U15010_Pad12, __A15_1__FB11, __A15_1__FB11_n, GND, net_U15010_Pad8, SUMA03_n, U2BBKG_n, SUMB03_n, net_U15010_Pad12, SUMB11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15011(net_U15011_Pad1, WL11_n, WEBG_n, net_U15011_Pad4, WL03_n, WBBEG_n, GND, EB11_n, CEBG, __A15_1__EB11, REBG_n, EB11_n, net_U15009_Pad12, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U15012(EB11_n, net_U15010_Pad8, net_U15011_Pad1, net_U15011_Pad4, __A15_1__EB11,  , GND,  , net_U15012_Pad9, net_U15012_Pad10, net_U15012_Pad11, EB10, __A15_1__EB10_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15013(__A15_1__BBK3, EB11_n, RBBEG_n, net_U15012_Pad10, WL10_n, WEBG_n, GND, WL02_n, WBBEG_n, net_U15012_Pad11, __A15_1__EB10_n, CEBG, EB10, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15014(SUMA02_n, U2BBKG_n, SUMA01_n, U2BBKG_n, SUMB01_n, net_U15014_Pad6, GND, __A15_1__F14, net_U15014_Pad9, net_U15014_Pad10, __A15_1__FB14_n, net_U15012_Pad9, SUMB02_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15015(net_U15003_Pad11, REBG_n, __A15_1__EB10_n, __A15_1__BBK2, __A15_1__EB10_n, RBBEG_n, GND, WL09_n, WEBG_n, net_U15015_Pad10, WL01_n, WBBEG_n, net_U15015_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15016(net_U15003_Pad10, RL10_n, net_U15003_Pad12, RL09_n, net_U15016_Pad5, RL06_n, GND, net_R15001_Pad2, net_U15016_Pad9, net_R15001_Pad2, net_U15016_Pad11, net_R15002_Pad2, net_U15016_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 #(1'b1, 1'b1) U15017(__A15_1__EB9_n, net_U15014_Pad6, net_U15015_Pad10, net_U15015_Pad13, EB9,  , GND,  , __A15_1__FB14_n, __A15_1__FB16_n, E7_n, net_U15014_Pad9, __A15_1__F16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15018(EB9, __A15_1__EB9_n, CEBG, net_U15003_Pad13, REBG_n, __A15_1__EB9_n, GND, __A15_1__EB9_n, RBBEG_n, __A15_1__BBK1, __A15_1__FB11_n, net_U15014_Pad9, net_U15018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15019(S12_n, net_U15014_Pad9, __A15_1__F11_n, __A15_1__F11, __A15_1__F12_n, __A15_1__F12, GND, __A15_1__F13_n, __A15_1__F13, __A15_1__F14_n, __A15_1__F14, __A15_1__F15_n, __A15_1__F15, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15020(__A15_1__F11_n, net_U15018_Pad13, net_U15020_Pad3, net_U15020_Pad3, S11_n, S12_n, GND, net_U15014_Pad9, __A15_1__FB12, __A15_1__F12_n, net_U15014_Pad9, __A15_1__FB13_n, __A15_1__F13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15021(E5, __A15_1__FB16_n, __A15_1__FB16_n, net_U15021_Pad4, net_U15014_Pad9, __A15_1__F15, GND, net_U15021_Pad4, E7_n, __A15_1__FB14_n, E6, net_U15014_Pad10, E7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15022(__A15_1__F16, __A15_1__F16_n, net_U15022_Pad3, net_U15022_Pad4, KRPT, __A15_1__KRPTA_n, GND, net_U15022_Pad8, net_U15022_Pad9, net_U15022_Pad10, net_U15022_Pad11, __A15_1__PRPOR1, net_U15022_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15023(XB4_n, XT4_n, __A15_1__KRPTA_n, XB0_n, XT5_n, net_U15023_Pad6, GND, net_U15023_Pad8, net_U15023_Pad9, net_U15023_Pad10, GOJAM, net_U15023_Pad10, __A15_1__KRPTA_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U15024(net_U15023_Pad9, RADRPT, net_U15023_Pad8, net_U15024_Pad4, HNDRPT, net_U15024_Pad6, GND, net_U15024_Pad8, __A15_1__RRPA1_n, __A15_1__RPTAD6, __A15_1__RRPA1_n, net_U15024_Pad12, __A15_1__RPTA12, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15025(net_U15024_Pad4, net_U15023_Pad6, __A15_1__PRPOR1, net_U15023_Pad9, __A15_1__DNRPTA, __A15_1__PRPOR3, GND, net_U15024_Pad8, __A15_1__PRPOR2, __A15_1__PRPOR3, __A15_1__PRPOR4, net_U15024_Pad6, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U15026(__A15_1__PRPOR4, __A15_1__PRPOR1, __A15_1__DNRPTA, net_U15023_Pad8, net_U15024_Pad4,  , GND,  , net_U15024_Pad6, net_U15023_Pad8, __A15_1__PRPOR1, __A15_1__DNRPTA, net_U15024_Pad12, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U15027(net_U15016_Pad5, CAD6, __A15_1__RPTAD6, net_U15027_Pad4, net_U15024_Pad12, RUPTOR_n, GND, net_U15027_Pad4, T10, RUPTOR_n, WOVR_n, OVF_n, net_U15022_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15028(CA3_n, XB1_n, net_U15028_Pad3, GOJAM, net_U15028_Pad5, net_U15028_Pad6, GND, net_U15028_Pad5, XT0_n, XB4_n, __A15_1__KRPTA_n, T6RPT, ZOUT_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U15029(net_U15028_Pad3, T6RPT, net_U15028_Pad6, net_U15029_Pad4, net_U15029_Pad5, net_U15029_Pad6, GND, net_U15029_Pad8, net_U15029_Pad9, net_U15029_Pad10, net_U15029_Pad11, net_U15029_Pad12, net_U15029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15030(CA3_n, XB0_n, net_U15029_Pad4, GOJAM, net_U15030_Pad5, net_U15029_Pad6, GND, net_U15030_Pad5, XB0_n, XT1_n, __A15_1__KRPTA_n, net_U15029_Pad5, net_U15022_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15031(CA2_n, XB6_n, net_U15029_Pad10, GOJAM, net_U15031_Pad5, net_U15029_Pad9, GND, net_U15031_Pad5, XT1_n, XB4_n, __A15_1__KRPTA_n, net_U15029_Pad8, net_U15022_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15032(CA2_n, XB7_n, net_U15029_Pad13, GOJAM, net_U15032_Pad5, net_U15029_Pad12, GND, net_U15032_Pad5, XT2_n, XB0_n, __A15_1__KRPTA_n, net_U15029_Pad11, net_U15022_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U15033(net_U15033_Pad1, KYRPT1, net_U15033_Pad3, net_U15033_Pad4, UPRUPT, net_U15033_Pad6, GND, DLKPLS, __A15_1__DNRPTA, net_U15033_Pad10, net_U15028_Pad6, net_U15029_Pad4, net_U15033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U15034(net_U15033_Pad1, GOJAM, XB4_n, XT2_n, __A15_1__KRPTA_n, __A15_2__KY1RST, GND, net_U15034_Pad8, KYRPT2, MKRPT, net_U15034_Pad11, net_U15033_Pad3, __A15_2__KY1RST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15035(net_U15034_Pad8, GOJAM, XT3_n, XB0_n, __A15_1__KRPTA_n, __A15_2__KY2RST, GND, net_U15033_Pad6, net_U15033_Pad4, GOJAM, net_U15035_Pad11, net_U15034_Pad11, __A15_2__KY2RST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15036(XT3_n, XB4_n, net_U15033_Pad10, GOJAM, DRPRST, __A15_1__DNRPTA, GND, DRPRST, XB0_n, XT4_n, __A15_1__KRPTA_n, net_U15035_Pad11, __A15_1__KRPTA_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15037(net_U15016_Pad9, net_U15028_Pad6, net_U15037_Pad3, net_U15016_Pad13, net_U15033_Pad13, net_U15037_Pad3, GND, net_U15022_Pad8, net_U15029_Pad13, net_U15037_Pad10, net_U15022_Pad10, net_U15034_Pad8, net_U15037_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15038(net_U15038_Pad1, net_U15038_Pad10, net_U15028_Pad6, net_U15029_Pad10, net_U15029_Pad6, net_U15037_Pad3, GND, net_U15038_Pad8, net_U15037_Pad13, net_U15038_Pad10, __A15_1__PRPOR4, net_U15016_Pad11, __A15_1__PRPOR3, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15039(net_U15038_Pad8, net_R15002_Pad2, net_U15039_Pad3, RL03_n, net_U15039_Pad5, RL04_n, GND, RL05_n, net_U15039_Pad9, RL02_n, net_U15039_Pad11, RL01_n, net_U15039_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U15040(net_U15028_Pad6, net_U15029_Pad9, net_U15022_Pad8, net_U15033_Pad1, net_U15029_Pad12, net_U15038_Pad1, GND, net_U15022_Pad11, net_U15022_Pad8, net_U15033_Pad3, net_U15029_Pad12, net_U15022_Pad9, net_U15029_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U15041(net_U15041_Pad1, net_U15038_Pad1, net_U15037_Pad10, net_U15037_Pad13, net_U15038_Pad10,  , GND,  , __A15_2__RPTAD3, __A15_1__BBK3, CAD3, R6, net_U15039_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15042(net_U15022_Pad10, net_U15033_Pad4, net_U15022_Pad10, net_U15033_Pad6, net_U15034_Pad11, net_U15022_Pad13, GND,  ,  ,  ,  , net_U15038_Pad10, net_U15034_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15043(__A15_1__PRPOR2, __A15_1__PRPOR1, net_U15033_Pad10, __A15_2__RPTAD3, __A15_1__RRPA1_n, net_R15001_Pad2, GND, __A15_1__RRPA1_n, net_R15002_Pad2, __A15_2__RPTAD4, __A15_2__RPTAD4, CAD4, net_U15039_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15044(RRPA, __A15_1__RRPA1_n, STRGAT, net_U15044_Pad4, __A15_1__F11, net_U15044_Pad6, GND, net_U15044_Pad8, __A15_1__F11_n, net_U15044_Pad10, S10, net_U15044_Pad12, S10_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15045(net_U15039_Pad9, __A15_2__RPTAD5, CAD5, __A15_2__RPTAD5, __A15_1__RRPA1_n, net_U15041_Pad1, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15046(CAD2, __A15_1__BBK2, CAD1, __A15_1__BBK1, RB1F, net_U15039_Pad13, GND, STR412, net_U15044_Pad4, net_U15044_Pad10, net_U15044_Pad6, net_U15039_Pad11, R6, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15047(net_U15044_Pad4, net_U15044_Pad12, net_U15044_Pad4, net_U15044_Pad10, net_U15044_Pad8, STR210, GND, STR19, net_U15044_Pad4, net_U15044_Pad12, net_U15044_Pad8, STR311, net_U15044_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15048(net_U15048_Pad1, __A15_1__F16, __A15_1__F15, net_U15048_Pad4, __A15_1__F16, __A15_1__F15_n, GND, __A15_1__F15, __A15_1__F16_n, net_U15048_Pad10, __A15_2__NE036_n, __A15_1__F12, __A15_2__036L, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15049(net_U15048_Pad1, net_U15049_Pad2, __A15_1__F14_n, net_U15049_Pad4, __A15_1__F13_n, net_U15049_Pad6, GND, net_U15049_Pad8, __A15_1__F13, net_U15049_Pad10, __A15_1__F14, net_U15049_Pad12, net_U15048_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15050(net_U15049_Pad2, net_U15049_Pad4, net_U15049_Pad2, net_U15049_Pad4, net_U15049_Pad8, __A15_2__NE01, GND, __A15_2__NE02, net_U15049_Pad2, net_U15049_Pad10, net_U15049_Pad6, __A15_2__NE00, net_U15049_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15051(net_U15049_Pad2, net_U15049_Pad10, net_U15049_Pad12, net_U15049_Pad4, net_U15049_Pad6, __A15_2__NE04, GND, __A15_2__NE05, net_U15049_Pad12, net_U15049_Pad4, net_U15049_Pad8, __A15_2__NE03, net_U15049_Pad8, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15052(net_U15049_Pad12, net_U15049_Pad10, net_U15049_Pad12, net_U15049_Pad10, net_U15049_Pad8, __A15_2__NE07, GND, __A15_2__NE10, net_U15052_Pad9, net_U15049_Pad4, net_U15049_Pad6, __A15_2__NE06, net_U15049_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15053(net_U15048_Pad10, net_U15052_Pad9, net_U15053_Pad3, STR14,  ,  , GND, LOMOD, net_U15053_Pad9, STR58, net_U15053_Pad11,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15054(__A15_2__NE00, __A15_2__NE03, __A15_2__NE00, __A15_2__NE01, __A15_2__NE02, __A15_2__NE012_n, GND, __A15_2__NE147_n, __A15_2__NE01, __A15_2__NE04, __A15_2__NE07, __A15_2__NE036_n, __A15_2__NE06, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15055(__A15_2__NE04, __A15_2__NE03, __A15_2__NE02, __A15_2__NE05, __A15_2__NE10, __A15_2__NE2510_n, GND, __A15_2__NE6710_n, __A15_2__NE06, __A15_2__NE07, __A15_2__NE10, __A15_2__NE345_n, __A15_2__NE05, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15056(__A15_2__147H, __A15_2__NE147_n, __A15_1__F12_n, __A15_2__2510L, __A15_2__NE2510_n, __A15_1__F12, GND, __A15_2__NE036_n, __A15_1__F12_n, __A15_2__036H, __A15_2__NE147_n, __A15_1__F12, __A15_2__147L, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15057(__A15_2__2510H, __A15_2__NE2510_n, __A15_1__F12_n, net_U15053_Pad3, __A15_2__036L, __A15_2__147H, GND, __A15_2__2510L, __A15_2__036H, net_U15053_Pad11, __A15_2__147L, __A15_2__2510H, net_U15057_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15058(__A15_2__036L, __A15_2__147L, __A15_2__147H, __A15_2__2510H, __A15_2__2510L, net_U15058_Pad6, GND,  ,  ,  ,  , net_U15053_Pad9, __A15_2__036H, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15059(net_U15058_Pad6, HIMOD, net_U15057_Pad13, STR912,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15060(ROPER, __A15_2__NE012_n, STRT2, ROPES, __A15_2__NE345_n, STRT2, GND, __A15_2__NE6710_n, STRT2, ROPET,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule