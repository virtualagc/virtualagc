`timescale 1ns/1ps
`default_nettype none

module inout_i(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, CCHG_n, WCHG_n, CCH11, RCH11_n, WCH11_n, FLASH, FLASH_n, XT0_n, XT1_n, XB2_n, XB5_n, XB6_n, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CH0705, CH0706, CH0707, CH1501, CH1502, CH1503, CH1504, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207, CH3208, CCH12, RCH12_n, WCH12_n, TMPOUT, CH1213, CH1214, CH1208, CH1209, CH1210, CH1211, CH1212, CHOR01_n, CHOR02_n, CHOR03_n, CHOR04_n, CHOR05_n, CHOR06_n, CHOR07_n, CHOR08_n, COMACT, UPLACT, KYRLS, VNFLSH, OPEROR);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire CCH11;
    output wire CCH12;
    input wire CCHG_n;
    input wire CH0705;
    input wire CH0706;
    input wire CH0707;
    output wire CH1208;
    output wire CH1209;
    output wire CH1210;
    output wire CH1211;
    output wire CH1212;
    output wire CH1213;
    output wire CH1214;
    input wire CH1501;
    input wire CH1502;
    input wire CH1503;
    input wire CH1504;
    input wire CH3201;
    input wire CH3202;
    input wire CH3203;
    input wire CH3204;
    input wire CH3205;
    input wire CH3206;
    input wire CH3207;
    input wire CH3208;
    output wire CHOR01_n; //FPGA#wand
    output wire CHOR02_n; //FPGA#wand
    output wire CHOR03_n; //FPGA#wand
    output wire CHOR04_n; //FPGA#wand
    output wire CHOR05_n; //FPGA#wand
    output wire CHOR06_n; //FPGA#wand
    output wire CHOR07_n; //FPGA#wand
    output wire CHOR08_n; //FPGA#wand
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    output wire COMACT;
    input wire FLASH;
    input wire FLASH_n;
    input wire GOJAM;
    output wire KYRLS;
    output wire OPEROR;
    input wire RCH11_n;
    output wire RCH12_n;
    output wire TMPOUT;
    output wire UPLACT;
    output wire VNFLSH;
    input wire WCH11_n;
    output wire WCH12_n;
    input wire WCHG_n;
    input wire XB2_n;
    input wire XB5_n;
    input wire XB6_n;
    input wire XT0_n;
    input wire XT1_n;
    wire __A16_1__CCH05;
    wire __A16_1__CCH06;
    wire __A16_1__CH1207;
    wire __A16_1__OT1207;
    wire __A16_1__OT1207_n;
    wire __A16_1__RCH05_n;
    wire __A16_1__RCH06_n;
    wire __A16_1__RCmXmP;
    wire __A16_1__RCmXmY;
    wire __A16_1__RCmXpP;
    wire __A16_1__RCmXpY;
    wire __A16_1__RCmYmR;
    wire __A16_1__RCmYpR;
    wire __A16_1__RCmZmR;
    wire __A16_1__RCmZpR;
    wire __A16_1__RCpXmP;
    wire __A16_1__RCpXmY;
    wire __A16_1__RCpXpP;
    wire __A16_1__RCpXpY;
    wire __A16_1__RCpYmR;
    wire __A16_1__RCpYpR;
    wire __A16_1__RCpZmR;
    wire __A16_1__RCpZpR;
    wire __A16_1__TVCNAB;
    wire __A16_1__WCH05_n;
    wire __A16_1__WCH06_n;
    wire __A16_2__COARSE;
    wire __A16_2__DISDAC;
    wire __A16_2__ENERIM;
    wire __A16_2__ENEROP;
    wire __A16_2__ISSWAR;
    wire __A16_2__MROLGT;
    wire __A16_2__S4BOFF;
    wire __A16_2__S4BSEQ;
    wire __A16_2__S4BTAK;
    wire __A16_2__STARON;
    wire __A16_2__ZEROPT;
    wire __A16_2__ZIMCDU;
    wire __A16_2__ZOPCDU;
    wire net_U16001_Pad1;
    wire net_U16001_Pad10;
    wire net_U16001_Pad11;
    wire net_U16001_Pad13;
    wire net_U16002_Pad11;
    wire net_U16002_Pad13;
    wire net_U16002_Pad3;
    wire net_U16002_Pad5;
    wire net_U16002_Pad9;
    wire net_U16003_Pad1;
    wire net_U16003_Pad10;
    wire net_U16003_Pad12;
    wire net_U16003_Pad3;
    wire net_U16003_Pad4;
    wire net_U16003_Pad6;
    wire net_U16003_Pad8;
    wire net_U16003_Pad9;
    wire net_U16004_Pad11;
    wire net_U16004_Pad13;
    wire net_U16004_Pad9;
    wire net_U16005_Pad1;
    wire net_U16005_Pad10;
    wire net_U16006_Pad1;
    wire net_U16006_Pad10;
    wire net_U16007_Pad1;
    wire net_U16007_Pad10;
    wire net_U16008_Pad1;
    wire net_U16008_Pad10;
    wire net_U16009_Pad1;
    wire net_U16009_Pad10;
    wire net_U16010_Pad1;
    wire net_U16010_Pad10;
    wire net_U16010_Pad11;
    wire net_U16010_Pad13;
    wire net_U16011_Pad11;
    wire net_U16011_Pad13;
    wire net_U16011_Pad3;
    wire net_U16011_Pad5;
    wire net_U16011_Pad9;
    wire net_U16012_Pad1;
    wire net_U16012_Pad10;
    wire net_U16012_Pad3;
    wire net_U16012_Pad4;
    wire net_U16012_Pad9;
    wire net_U16013_Pad1;
    wire net_U16013_Pad10;
    wire net_U16014_Pad1;
    wire net_U16014_Pad10;
    wire net_U16015_Pad1;
    wire net_U16015_Pad10;
    wire net_U16016_Pad1;
    wire net_U16016_Pad10;
    wire net_U16017_Pad1;
    wire net_U16017_Pad10;
    wire net_U16018_Pad1;
    wire net_U16018_Pad10;
    wire net_U16018_Pad11;
    wire net_U16018_Pad13;
    wire net_U16019_Pad11;
    wire net_U16019_Pad13;
    wire net_U16019_Pad3;
    wire net_U16019_Pad5;
    wire net_U16019_Pad9;
    wire net_U16020_Pad1;
    wire net_U16020_Pad12;
    wire net_U16020_Pad3;
    wire net_U16020_Pad4;
    wire net_U16020_Pad6;
    wire net_U16021_Pad11;
    wire net_U16021_Pad13;
    wire net_U16021_Pad5;
    wire net_U16021_Pad9;
    wire net_U16022_Pad1;
    wire net_U16022_Pad10;
    wire net_U16023_Pad1;
    wire net_U16023_Pad10;
    wire net_U16024_Pad1;
    wire net_U16024_Pad10;
    wire net_U16025_Pad6;
    wire net_U16025_Pad8;
    wire net_U16026_Pad1;
    wire net_U16026_Pad11;
    wire net_U16026_Pad13;
    wire net_U16026_Pad3;
    wire net_U16026_Pad5;
    wire net_U16026_Pad9;
    wire net_U16028_Pad1;
    wire net_U16028_Pad10;
    wire net_U16029_Pad1;
    wire net_U16029_Pad10;
    wire net_U16030_Pad11;
    wire net_U16030_Pad13;
    wire net_U16030_Pad3;
    wire net_U16030_Pad5;
    wire net_U16030_Pad9;
    wire net_U16031_Pad1;
    wire net_U16031_Pad10;
    wire net_U16031_Pad13;
    wire net_U16032_Pad10;
    wire net_U16032_Pad2;
    wire net_U16032_Pad3;
    wire net_U16032_Pad4;
    wire net_U16032_Pad9;
    wire net_U16033_Pad1;
    wire net_U16033_Pad10;
    wire net_U16034_Pad1;
    wire net_U16034_Pad10;
    wire net_U16035_Pad1;
    wire net_U16035_Pad10;
    wire net_U16036_Pad1;
    wire net_U16036_Pad10;
    wire net_U16037_Pad1;
    wire net_U16037_Pad10;
    wire net_U16037_Pad11;
    wire net_U16038_Pad11;
    wire net_U16038_Pad13;
    wire net_U16038_Pad3;
    wire net_U16038_Pad5;
    wire net_U16038_Pad9;
    wire net_U16039_Pad1;
    wire net_U16039_Pad10;
    wire net_U16039_Pad13;
    wire net_U16040_Pad1;
    wire net_U16040_Pad10;
    wire net_U16040_Pad13;
    wire net_U16041_Pad10;
    wire net_U16041_Pad3;
    wire net_U16041_Pad4;
    wire net_U16041_Pad6;
    wire net_U16041_Pad8;
    wire net_U16041_Pad9;
    wire net_U16042_Pad1;
    wire net_U16042_Pad10;
    wire net_U16043_Pad1;
    wire net_U16043_Pad10;
    wire net_U16043_Pad11;
    wire net_U16044_Pad5;
    wire net_U16045_Pad1;
    wire net_U16045_Pad10;
    wire net_U16046_Pad1;
    wire net_U16046_Pad10;
    wire net_U16046_Pad11;
    wire net_U16047_Pad11;
    wire net_U16047_Pad13;
    wire net_U16047_Pad8;
    wire net_U16048_Pad1;
    wire net_U16048_Pad10;
    wire net_U16049_Pad1;
    wire net_U16049_Pad10;
    wire net_U16049_Pad11;
    wire net_U16050_Pad11;
    wire net_U16050_Pad13;
    wire net_U16050_Pad3;
    wire net_U16050_Pad5;
    wire net_U16050_Pad9;
    wire net_U16051_Pad1;
    wire net_U16051_Pad10;
    wire net_U16052_Pad1;
    wire net_U16052_Pad10;
    wire net_U16052_Pad13;
    wire net_U16054_Pad1;
    wire net_U16054_Pad10;
    wire net_U16055_Pad1;
    wire net_U16055_Pad10;
    wire net_U16056_Pad1;
    wire net_U16056_Pad10;
    wire net_U16057_Pad3;

    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16001(net_U16001_Pad1, CHWL01_n, __A16_1__WCH05_n, net_U16001_Pad11, net_U16001_Pad1, net_U16001_Pad10, GND, net_U16001_Pad11, __A16_1__CCH05, net_U16001_Pad10, net_U16001_Pad11, __A16_1__RCH05_n, net_U16001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16002(net_U16001_Pad11, __A16_1__RCpXpP, net_U16002_Pad3, __A16_1__RCpZpR, net_U16002_Pad5, __A16_1__RCmXmP, GND, __A16_1__RCmZmR, net_U16002_Pad9, __A16_1__RCmXpP, net_U16002_Pad11, __A16_1__RCmZpR, net_U16002_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16003(net_U16003_Pad1, net_U16001_Pad13, net_U16003_Pad3, net_U16003_Pad4, CH3202, net_U16003_Pad6, GND, net_U16003_Pad8, net_U16003_Pad9, net_U16003_Pad10, CH3203, net_U16003_Pad12, CH3201, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U16004(net_U16003_Pad12, CHOR01_n, net_U16003_Pad6, CHOR02_n, net_U16003_Pad8, CHOR03_n, GND, CHOR04_n, net_U16004_Pad9, CHOR05_n, net_U16004_Pad11, CHOR06_n, net_U16004_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16005(net_U16005_Pad1, CHWL01_n, __A16_1__WCH06_n, net_U16002_Pad3, net_U16005_Pad1, net_U16005_Pad10, GND, net_U16002_Pad3, __A16_1__CCH06, net_U16005_Pad10, net_U16002_Pad3, __A16_1__RCH06_n, net_U16003_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16006(net_U16006_Pad1, CHWL02_n, __A16_1__WCH05_n, net_U16002_Pad5, net_U16006_Pad1, net_U16006_Pad10, GND, net_U16002_Pad5, __A16_1__CCH05, net_U16006_Pad10, net_U16002_Pad5, __A16_1__RCH05_n, net_U16003_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16007(net_U16007_Pad1, CHWL02_n, __A16_1__WCH06_n, net_U16002_Pad9, net_U16007_Pad1, net_U16007_Pad10, GND, net_U16002_Pad9, __A16_1__CCH06, net_U16007_Pad10, net_U16002_Pad9, __A16_1__RCH06_n, net_U16003_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16008(net_U16008_Pad1, CHWL03_n, __A16_1__WCH05_n, net_U16002_Pad11, net_U16008_Pad1, net_U16008_Pad10, GND, net_U16002_Pad11, __A16_1__CCH05, net_U16008_Pad10, net_U16002_Pad11, __A16_1__RCH05_n, net_U16003_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16009(net_U16009_Pad1, CHWL03_n, __A16_1__WCH06_n, net_U16002_Pad13, net_U16009_Pad1, net_U16009_Pad10, GND, net_U16002_Pad13, __A16_1__CCH06, net_U16009_Pad10, net_U16002_Pad13, __A16_1__RCH06_n, net_U16003_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16010(net_U16010_Pad1, CHWL04_n, __A16_1__WCH05_n, net_U16010_Pad11, net_U16010_Pad1, net_U16010_Pad10, GND, net_U16010_Pad11, __A16_1__CCH05, net_U16010_Pad10, net_U16010_Pad11, __A16_1__RCH05_n, net_U16010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16011(net_U16010_Pad11, __A16_1__RCpXmP, net_U16011_Pad3, __A16_1__RCpZmR, net_U16011_Pad5, __A16_1__RCpXpY, GND, __A16_1__RCpYpR, net_U16011_Pad9, __A16_1__RCmXmY, net_U16011_Pad11, __A16_1__RCmYmR, net_U16011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16012(net_U16012_Pad1, net_U16010_Pad13, net_U16012_Pad3, net_U16012_Pad4, CH3205, net_U16004_Pad11, GND, net_U16004_Pad13, net_U16012_Pad9, net_U16012_Pad10, CH3206, net_U16004_Pad9, CH3204, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16013(net_U16013_Pad1, CHWL04_n, __A16_1__WCH06_n, net_U16011_Pad3, net_U16013_Pad1, net_U16013_Pad10, GND, net_U16011_Pad3, __A16_1__CCH06, net_U16013_Pad10, net_U16011_Pad3, __A16_1__RCH06_n, net_U16012_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16014(net_U16014_Pad1, CHWL05_n, __A16_1__WCH05_n, net_U16011_Pad5, net_U16014_Pad1, net_U16014_Pad10, GND, net_U16011_Pad5, __A16_1__CCH05, net_U16014_Pad10, net_U16011_Pad5, __A16_1__RCH05_n, net_U16012_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16015(net_U16015_Pad1, CHWL05_n, __A16_1__WCH06_n, net_U16011_Pad9, net_U16015_Pad1, net_U16015_Pad10, GND, net_U16011_Pad9, __A16_1__CCH06, net_U16015_Pad10, net_U16011_Pad9, __A16_1__RCH06_n, net_U16012_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16016(net_U16016_Pad1, CHWL06_n, __A16_1__WCH05_n, net_U16011_Pad11, net_U16016_Pad1, net_U16016_Pad10, GND, net_U16011_Pad11, __A16_1__CCH05, net_U16016_Pad10, net_U16011_Pad11, __A16_1__RCH05_n, net_U16012_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16017(net_U16017_Pad1, CHWL06_n, __A16_1__WCH06_n, net_U16011_Pad13, net_U16017_Pad1, net_U16017_Pad10, GND, net_U16011_Pad13, __A16_1__CCH06, net_U16017_Pad10, net_U16011_Pad13, __A16_1__RCH06_n, net_U16012_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16018(net_U16018_Pad1, CHWL07_n, __A16_1__WCH05_n, net_U16018_Pad11, net_U16018_Pad1, net_U16018_Pad10, GND, net_U16018_Pad11, __A16_1__CCH05, net_U16018_Pad10, net_U16018_Pad11, __A16_1__RCH05_n, net_U16018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16019(net_U16018_Pad11, __A16_1__RCmXpY, net_U16019_Pad3, __A16_1__RCmYpR, net_U16019_Pad5, __A16_1__RCpXmY, GND, __A16_1__RCpYmR, net_U16019_Pad9, __A16_1__WCH05_n, net_U16019_Pad11, __A16_1__WCH06_n, net_U16019_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16020(net_U16020_Pad1, net_U16018_Pad13, net_U16020_Pad3, net_U16020_Pad4, CH3208, net_U16020_Pad6, GND, net_U16019_Pad11, WCHG_n, XT0_n, XB5_n, net_U16020_Pad12, CH3207, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U16021(net_U16020_Pad12, CHOR07_n, net_U16020_Pad6, CHOR08_n, net_U16021_Pad5, CHOR01_n, GND, CHOR02_n, net_U16021_Pad9, CHOR03_n, net_U16021_Pad11, CHOR04_n, net_U16021_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16022(net_U16022_Pad1, CHWL07_n, __A16_1__WCH06_n, net_U16019_Pad3, net_U16022_Pad1, net_U16022_Pad10, GND, net_U16019_Pad3, __A16_1__CCH06, net_U16022_Pad10, net_U16019_Pad3, __A16_1__RCH06_n, net_U16020_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16023(net_U16023_Pad1, CHWL08_n, __A16_1__WCH05_n, net_U16019_Pad5, net_U16023_Pad1, net_U16023_Pad10, GND, net_U16019_Pad5, __A16_1__CCH05, net_U16023_Pad10, net_U16019_Pad5, __A16_1__RCH05_n, net_U16020_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16024(net_U16024_Pad1, CHWL08_n, __A16_1__WCH06_n, net_U16019_Pad9, net_U16024_Pad1, net_U16024_Pad10, GND, net_U16019_Pad9, __A16_1__CCH06, net_U16024_Pad10, net_U16019_Pad9, __A16_1__RCH06_n, net_U16020_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16025(WCHG_n, XT0_n, CCHG_n, XT0_n, XB5_n, net_U16025_Pad6, GND, net_U16025_Pad8, CCHG_n, XT0_n, XB6_n, net_U16019_Pad13, XB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16026(net_U16026_Pad1, __A16_1__CCH05, net_U16026_Pad3, __A16_1__RCH05_n, net_U16026_Pad5, __A16_1__RCH06_n, GND, __A16_1__CCH06, net_U16026_Pad9, __A16_1__TVCNAB, net_U16026_Pad11, __A16_1__OT1207, net_U16026_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U16027(net_U16026_Pad1, net_U16025_Pad6, GOJAM, net_U16026_Pad3, XT0_n, XB5_n, GND, XT0_n, XB6_n, net_U16026_Pad5, net_U16025_Pad8, GOJAM, net_U16026_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16028(net_U16028_Pad1, CHWL08_n, WCH12_n, net_U16026_Pad11, net_U16028_Pad1, net_U16028_Pad10, GND, net_U16026_Pad11, CCH12, net_U16028_Pad10, RCH12_n, net_U16026_Pad11, CH1208, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16029(net_U16029_Pad1, WCH12_n, CHWL07_n, net_U16026_Pad13, net_U16029_Pad1, net_U16029_Pad10, GND, net_U16026_Pad13, CCH12, net_U16029_Pad10, RCH12_n, net_U16026_Pad13, __A16_1__CH1207, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16030(net_U16029_Pad10, __A16_1__OT1207_n, net_U16030_Pad3, __A16_2__ZOPCDU, net_U16030_Pad5, __A16_2__ISSWAR, GND, __A16_2__ENEROP, net_U16030_Pad9, COMACT, net_U16030_Pad11, __A16_2__STARON, net_U16030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16031(net_U16031_Pad1, CHWL01_n, WCH12_n, net_U16030_Pad3, net_U16031_Pad1, net_U16031_Pad10, GND, net_U16030_Pad3, CCH12, net_U16031_Pad10, net_U16030_Pad3, RCH12_n, net_U16031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16032(net_U16031_Pad13, net_U16032_Pad2, net_U16032_Pad3, net_U16032_Pad4, CH1502, net_U16021_Pad9, GND, net_U16021_Pad11, net_U16032_Pad9, net_U16032_Pad10, CH1503, net_U16021_Pad5, CH1501, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16033(net_U16033_Pad1, CHWL01_n, WCH11_n, net_U16030_Pad5, net_U16033_Pad1, net_U16033_Pad10, GND, net_U16030_Pad5, CCH11, net_U16033_Pad10, net_U16030_Pad5, RCH11_n, net_U16032_Pad2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16034(net_U16034_Pad1, CHWL02_n, WCH12_n, net_U16030_Pad9, net_U16034_Pad1, net_U16034_Pad10, GND, net_U16030_Pad9, CCH12, net_U16034_Pad10, net_U16030_Pad9, RCH12_n, net_U16032_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16035(net_U16035_Pad1, CHWL02_n, WCH11_n, net_U16030_Pad11, net_U16035_Pad1, net_U16035_Pad10, GND, net_U16030_Pad11, CCH11, net_U16035_Pad10, net_U16030_Pad11, RCH11_n, net_U16032_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16036(net_U16036_Pad1, CHWL03_n, WCH12_n, net_U16030_Pad13, net_U16036_Pad1, net_U16036_Pad10, GND, net_U16030_Pad13, CCH12, net_U16036_Pad10, net_U16030_Pad13, RCH12_n, net_U16032_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16037(net_U16037_Pad1, CHWL03_n, WCH11_n, net_U16037_Pad11, net_U16037_Pad1, net_U16037_Pad10, GND, net_U16037_Pad11, CCH11, net_U16037_Pad10, net_U16037_Pad11, RCH11_n, net_U16032_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16038(net_U16037_Pad11, UPLACT, net_U16038_Pad3, __A16_2__COARSE, net_U16038_Pad5, TMPOUT, GND, __A16_2__ZIMCDU, net_U16038_Pad9, __A16_2__ENERIM, net_U16038_Pad11, __A16_2__S4BTAK, net_U16038_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16039(net_U16039_Pad1, CHWL04_n, WCH12_n, net_U16038_Pad3, net_U16039_Pad1, net_U16039_Pad10, GND, net_U16038_Pad3, CCH12, net_U16039_Pad10, net_U16038_Pad3, RCH12_n, net_U16039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16040(net_U16040_Pad1, CHWL04_n, WCH11_n, net_U16038_Pad5, net_U16040_Pad1, net_U16040_Pad10, GND, net_U16038_Pad5, CCH11, net_U16040_Pad10, net_U16038_Pad5, RCH11_n, net_U16040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16041(net_U16039_Pad13, net_U16040_Pad13, net_U16041_Pad3, net_U16041_Pad4, CH0705, net_U16041_Pad6, GND, net_U16041_Pad8, net_U16041_Pad9, net_U16041_Pad10, CH0706, net_U16021_Pad13, CH1504, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16042(net_U16042_Pad1, CHWL05_n, WCH12_n, net_U16038_Pad9, net_U16042_Pad1, net_U16042_Pad10, GND, net_U16038_Pad9, CCH12, net_U16042_Pad10, net_U16038_Pad9, RCH12_n, net_U16041_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16043(net_U16043_Pad1, CHWL05_n, WCH11_n, net_U16043_Pad11, net_U16043_Pad1, net_U16043_Pad10, GND, net_U16043_Pad11, CCH11, net_U16043_Pad10, net_U16043_Pad11, RCH11_n, net_U16041_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U16044(net_U16041_Pad6, CHOR05_n, net_U16041_Pad8, CHOR06_n, net_U16044_Pad5, CHOR07_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16045(net_U16045_Pad1, CHWL06_n, WCH12_n, net_U16038_Pad11, net_U16045_Pad1, net_U16045_Pad10, GND, net_U16038_Pad11, CCH12, net_U16045_Pad10, net_U16038_Pad11, RCH12_n, net_U16041_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16046(net_U16046_Pad1, CHWL06_n, WCH11_n, net_U16046_Pad11, net_U16046_Pad1, net_U16046_Pad10, GND, net_U16046_Pad11, CCH11, net_U16046_Pad10, net_U16046_Pad11, RCH11_n, net_U16041_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U16047(KYRLS, net_U16043_Pad11, FLASH, VNFLSH, net_U16046_Pad11, FLASH_n, GND, net_U16047_Pad8, FLASH, OPEROR, net_U16047_Pad11, GOJAM, net_U16047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16048(net_U16048_Pad1, CHWL09_n, WCH12_n, net_U16038_Pad13, net_U16048_Pad1, net_U16048_Pad10, GND, net_U16038_Pad13, CCH12, net_U16048_Pad10, net_U16038_Pad13, RCH12_n, CH1209, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16049(net_U16049_Pad1, CHWL10_n, WCH12_n, net_U16049_Pad11, net_U16049_Pad1, net_U16049_Pad10, GND, net_U16049_Pad11, CCH12, net_U16049_Pad10, net_U16049_Pad11, RCH12_n, CH1210, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16050(net_U16049_Pad11, __A16_2__ZEROPT, net_U16050_Pad3, __A16_2__DISDAC, net_U16050_Pad5, __A16_2__MROLGT, GND, __A16_2__S4BSEQ, net_U16050_Pad9, __A16_2__S4BOFF, net_U16050_Pad11, WCH12_n, net_U16050_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16051(net_U16051_Pad1, CHWL11_n, WCH12_n, net_U16050_Pad3, net_U16051_Pad1, net_U16051_Pad10, GND, net_U16050_Pad3, CCH12, net_U16051_Pad10, net_U16050_Pad3, RCH12_n, CH1211, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16052(net_U16052_Pad1, CHWL07_n, WCH11_n, net_U16047_Pad8, net_U16052_Pad1, net_U16052_Pad10, GND, net_U16047_Pad8, CCH11, net_U16052_Pad10, net_U16047_Pad8, RCH11_n, net_U16052_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16053(__A16_1__CH1207, net_U16052_Pad13, WCHG_n, XB2_n, XT1_n, net_U16050_Pad13, GND, net_U16047_Pad11, CCHG_n, XB2_n, XT1_n, net_U16044_Pad5, CH0707, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16054(net_U16054_Pad1, CHWL12_n, WCH12_n, net_U16050_Pad5, net_U16054_Pad1, net_U16054_Pad10, GND, net_U16050_Pad5, CCH12, net_U16054_Pad10, net_U16050_Pad5, RCH12_n, CH1212, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16055(net_U16055_Pad1, CHWL13_n, WCH12_n, net_U16050_Pad9, net_U16055_Pad1, net_U16055_Pad10, GND, net_U16050_Pad9, CCH12, net_U16055_Pad10, net_U16050_Pad9, RCH12_n, CH1213, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16056(net_U16056_Pad1, CHWL14_n, WCH12_n, net_U16050_Pad11, net_U16056_Pad1, net_U16056_Pad10, GND, net_U16050_Pad11, CCH12, net_U16056_Pad10, net_U16050_Pad11, RCH12_n, CH1214, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16057(net_U16047_Pad13, CCH12, net_U16057_Pad3, RCH12_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U16058(net_U16057_Pad3, XT1_n, XB2_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule