`timescale 1ns/1ps
`default_nettype none

module counter_cell_ii(SIM_RST, SIM_CLK, p4VSW, GND, T12, T12A, INCSET_n, RSCT, BKTF_n, RSSB, BMAGXP, BMAGXM, BMAGYP, BMAGYM, EMSD, OTLNKM, ALTM, BMAGZP, BMAGZM, INLNKP, INLNKM, RNRADP, RNRADM, GYROD, XB0, XB1, XB2, XB3, XB4, XB5, XB6, XB7, OCTAD2, OCTAD3, OCTAD4, OCTAD5, OCTAD6, CG13, CG23, C24A, C25A, C26A, C27A, C30A, C31A, C32A, C32P, C32M, C33A, C33P, C33M, C34A, C34P, C34M, C35A, C35P, C35M, C36A, C36P, C36M, C37A, C37P, C37M, C40A, C40P, C40M, C41A, C41P, C41M, C50A, C51A, C52A, C53A, C54A, C55A, CA2_n, CA3_n, CA4_n, CA5_n, CA6_n, CXB0_n, CXB1_n, CXB2_n, CXB3_n, CXB4_n, CXB5_n, CXB6_n, CXB7_n, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CG26, C45R, PINC, MINC, DINC, DINC_n, PCDU, MCDU, SHINC_n, SHANC_n, SHIFT, SHIFT_n, CTROR, CTROR_n);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire ALTM;
    input wire BKTF_n;
    input wire BMAGXM;
    input wire BMAGXP;
    input wire BMAGYM;
    input wire BMAGYP;
    input wire BMAGZM;
    input wire BMAGZP;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C31A;
    input wire C32A;
    input wire C32M;
    input wire C32P;
    input wire C33A;
    input wire C33M;
    input wire C33P;
    input wire C34A;
    input wire C34M;
    input wire C34P;
    input wire C35A;
    input wire C35M;
    input wire C35P;
    input wire C36A;
    input wire C36M;
    input wire C36P;
    input wire C37A;
    input wire C37M;
    input wire C37P;
    input wire C40A;
    input wire C40M;
    input wire C40P;
    input wire C41A;
    input wire C41M;
    input wire C41P;
    output wire C45R;
    input wire C50A;
    input wire C51A;
    input wire C52A;
    input wire C53A;
    input wire C54A;
    input wire C55A;
    output wire CA2_n;
    output wire CA3_n;
    output wire CA4_n;
    output wire CA5_n;
    output wire CA6_n;
    output wire CAD1;
    output wire CAD2;
    output wire CAD3;
    output wire CAD4;
    output wire CAD5;
    output wire CAD6;
    input wire CG13;
    input wire CG23;
    output wire CG26;
    output wire CTROR;
    output wire CTROR_n;
    output wire CXB0_n;
    output wire CXB1_n;
    output wire CXB2_n;
    output wire CXB3_n;
    output wire CXB4_n;
    output wire CXB5_n;
    output wire CXB6_n;
    output wire CXB7_n;
    output wire DINC;
    output wire DINC_n;
    input wire EMSD;
    input wire GYROD;
    input wire INCSET_n;
    input wire INLNKM;
    input wire INLNKP;
    output wire MCDU;
    output wire MINC;
    input wire OCTAD2;
    input wire OCTAD3;
    input wire OCTAD4;
    input wire OCTAD5;
    input wire OCTAD6;
    input wire OTLNKM;
    output wire PCDU;
    output wire PINC;
    input wire RNRADM;
    input wire RNRADP;
    input wire RSCT;
    input wire RSSB;
    output wire SHANC_n;
    output wire SHIFT;
    output wire SHIFT_n;
    output wire SHINC_n;
    input wire T12;
    input wire T12A;
    input wire XB0;
    input wire XB1;
    input wire XB2;
    input wire XB3;
    input wire XB4;
    input wire XB5;
    input wire XB6;
    input wire XB7;
    wire __A21_1__30SUM;
    wire __A21_1__32004K; //FPGA#wand
    wire __A21_1__50SUM;
    wire __A21_1__C42A;
    wire __A21_1__C42M;
    wire __A21_1__C42P;
    wire __A21_1__C43A;
    wire __A21_1__C43M;
    wire __A21_1__C43P;
    wire __A21_1__C44A;
    wire __A21_1__C44M;
    wire __A21_1__C44P;
    wire __A21_1__C45A;
    wire __A21_1__C45M;
    wire __A21_1__C45P;
    wire __A21_1__C46A;
    wire __A21_1__C46M;
    wire __A21_1__C46P;
    wire __A21_1__C47A;
    wire __A21_1__C56A;
    wire __A21_1__C57A;
    wire __A21_1__C60A;
    wire __A21_1__DINCNC_n;
    wire __A21_1__MCDU_n;
    wire __A21_1__MINC_n;
    wire __A21_1__PCDU_n;
    wire __A21_1__PINC_n;
    wire __A21_1__RSCT_n;
    wire __A21_1__SHANC;
    wire __A21_1__SHINC;
    wire __A21_3__C42R;
    wire __A21_3__C43R;
    wire __A21_3__C44R;
    wire __A21_3__C46R;
    wire __A21_3__C47R;
    wire __A21_3__C56R;
    wire __A21_3__C57R;
    wire __A21_3__C60R;
    wire __A21_3__CG15;
    wire __A21_3__CG16;
    wire net_R21001_Pad2; //FPGA#wand
    wire net_R21002_Pad2; //FPGA#wand
    wire net_R21003_Pad2; //FPGA#wand
    wire net_R21005_Pad2; //FPGA#wand
    wire net_R21006_Pad2; //FPGA#wand
    wire net_R21007_Pad2; //FPGA#wand
    wire net_R21008_Pad2; //FPGA#wand
    wire net_R21009_Pad2; //FPGA#wand
    wire net_R21010_Pad2; //FPGA#wand
    wire net_R21011_Pad2; //FPGA#wand
    wire net_R21012_Pad2; //FPGA#wand
    wire net_U21001_Pad1;
    wire net_U21001_Pad13;
    wire net_U21002_Pad11;
    wire net_U21002_Pad13;
    wire net_U21002_Pad5;
    wire net_U21002_Pad9;
    wire net_U21004_Pad10;
    wire net_U21004_Pad13;
    wire net_U21004_Pad4;
    wire net_U21005_Pad13;
    wire net_U21006_Pad11;
    wire net_U21006_Pad13;
    wire net_U21006_Pad5;
    wire net_U21006_Pad9;
    wire net_U21009_Pad1;
    wire net_U21009_Pad13;
    wire net_U21010_Pad11;
    wire net_U21010_Pad5;
    wire net_U21010_Pad9;
    wire net_U21013_Pad13;
    wire net_U21014_Pad11;
    wire net_U21014_Pad13;
    wire net_U21014_Pad3;
    wire net_U21014_Pad9;
    wire net_U21015_Pad13;
    wire net_U21016_Pad1;
    wire net_U21017_Pad13;
    wire net_U21019_Pad1;
    wire net_U21019_Pad10;
    wire net_U21019_Pad4;
    wire net_U21021_Pad4;
    wire net_U21022_Pad1;
    wire net_U21022_Pad13;
    wire net_U21023_Pad11;
    wire net_U21023_Pad13;
    wire net_U21023_Pad5;
    wire net_U21023_Pad9;
    wire net_U21025_Pad1;
    wire net_U21025_Pad13;
    wire net_U21026_Pad6;
    wire net_U21027_Pad5;
    wire net_U21028_Pad1;
    wire net_U21029_Pad1;
    wire net_U21029_Pad11;
    wire net_U21029_Pad13;
    wire net_U21030_Pad1;
    wire net_U21030_Pad10;
    wire net_U21030_Pad13;
    wire net_U21030_Pad3;
    wire net_U21031_Pad10;
    wire net_U21031_Pad12;
    wire net_U21031_Pad2;
    wire net_U21031_Pad4;
    wire net_U21031_Pad5;
    wire net_U21032_Pad1;
    wire net_U21032_Pad10;
    wire net_U21032_Pad13;
    wire net_U21032_Pad4;
    wire net_U21033_Pad12;
    wire net_U21033_Pad13;
    wire net_U21035_Pad10;
    wire net_U21035_Pad12;
    wire net_U21035_Pad13;
    wire net_U21035_Pad4;
    wire net_U21036_Pad10;
    wire net_U21036_Pad12;
    wire net_U21036_Pad13;
    wire net_U21039_Pad1;
    wire net_U21039_Pad12;
    wire net_U21039_Pad13;
    wire net_U21039_Pad3;
    wire net_U21040_Pad10;
    wire net_U21040_Pad13;
    wire net_U21040_Pad4;
    wire net_U21042_Pad1;
    wire net_U21042_Pad10;
    wire net_U21042_Pad12;
    wire net_U21042_Pad13;
    wire net_U21042_Pad3;
    wire net_U21043_Pad10;
    wire net_U21043_Pad12;
    wire net_U21043_Pad13;
    wire net_U21043_Pad4;
    wire net_U21045_Pad10;
    wire net_U21045_Pad12;
    wire net_U21045_Pad13;
    wire net_U21045_Pad4;
    wire net_U21045_Pad7;
    wire net_U21046_Pad10;
    wire net_U21046_Pad13;
    wire net_U21048_Pad1;
    wire net_U21048_Pad10;
    wire net_U21048_Pad13;
    wire net_U21048_Pad3;
    wire net_U21049_Pad1;
    wire net_U21049_Pad10;
    wire net_U21049_Pad13;
    wire net_U21049_Pad3;
    wire net_U21051_Pad6;
    wire net_U21052_Pad3;
    wire net_U21053_Pad1;
    wire net_U21053_Pad10;
    wire net_U21053_Pad12;
    wire net_U21053_Pad3;
    wire net_U21054_Pad1;
    wire net_U21054_Pad11;
    wire net_U21054_Pad12;
    wire net_U21054_Pad13;
    wire net_U21054_Pad3;
    wire net_U21055_Pad10;
    wire net_U21055_Pad12;

    pullup R21001(net_R21001_Pad2);
    pullup R21002(net_R21002_Pad2);
    pullup R21003(net_R21003_Pad2);
    pullup R21004(__A21_1__32004K);
    pullup R21005(net_R21005_Pad2);
    pullup R21006(net_R21006_Pad2);
    pullup R21007(net_R21007_Pad2);
    pullup R21008(net_R21008_Pad2);
    pullup R21009(net_R21009_Pad2);
    pullup R21010(net_R21010_Pad2);
    pullup R21011(net_R21011_Pad2);
    pullup R21012(net_R21012_Pad2);
    U74HC4002 U21001(net_U21001_Pad1, C25A, C27A, C31A, C33A,  , GND,  , C35A, C37A, C41A, __A21_1__C43A, net_U21001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21002(net_U21001_Pad1, net_R21001_Pad2, net_U21001_Pad13, net_R21001_Pad2, net_U21002_Pad5, net_R21001_Pad2, GND, net_R21001_Pad2, net_U21002_Pad9, net_R21002_Pad2, net_U21002_Pad11, net_R21002_Pad2, net_U21002_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21003(net_U21002_Pad5, __A21_1__C45A, __A21_1__C47A, C51A, C53A,  , GND,  , C26A, C27A, C32A, C33A, net_U21002_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21004(net_U21002_Pad9, C55A, __A21_1__C57A, net_U21004_Pad4, __A21_1__C56A, __A21_1__C57A, GND, __A21_1__30SUM, __A21_1__C60A, net_U21004_Pad10, __A21_1__50SUM, __A21_1__C60A, net_U21004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21005(net_U21002_Pad13, C36A, C37A, __A21_1__C42A, __A21_1__C43A,  , GND,  , __A21_1__C46A, __A21_1__C47A, C52A, C53A, net_U21005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21006(net_U21005_Pad13, net_R21002_Pad2, net_U21004_Pad4, net_R21002_Pad2, net_U21006_Pad5, net_R21003_Pad2, GND, net_R21003_Pad2, net_U21006_Pad9, net_R21003_Pad2, net_U21006_Pad11, net_R21003_Pad2, net_U21006_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21007(net_U21006_Pad5, C24A, C25A, C26A, C27A,  , GND,  , C34A, C35A, C36A, C37A, net_U21006_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21008(net_U21006_Pad11, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, net_U21006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21009(net_U21009_Pad1, C30A, C31A, C32A, C33A,  , GND,  , C34A, C35A, C36A, C37A, net_U21009_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21010(net_U21009_Pad1, __A21_1__32004K, net_U21009_Pad13, __A21_1__32004K, net_U21010_Pad5, net_R21005_Pad2, GND, net_R21005_Pad2, net_U21010_Pad9, net_R21006_Pad2, net_U21010_Pad11, net_R21006_Pad2, net_U21004_Pad10, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC04 U21011(__A21_1__32004K, __A21_1__30SUM, net_R21005_Pad2, __A21_1__50SUM, DINC, DINC_n, GND, CXB0_n, XB0, CXB1_n, XB1, CXB2_n, XB2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21012(net_U21010_Pad5, C50A, C51A, C52A, C53A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, net_U21010_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21013(net_U21010_Pad11, C24A, C25A, C26A, C27A,  , GND,  , C40A, C41A, __A21_1__C42A, __A21_1__C43A, net_U21013_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21014(net_U21013_Pad13, net_R21007_Pad2, net_U21014_Pad3, net_R21007_Pad2, net_U21004_Pad13, net_R21007_Pad2, GND, net_R21008_Pad2, net_U21014_Pad9, net_R21008_Pad2, net_U21014_Pad11, net_R21008_Pad2, net_U21014_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21015(net_U21014_Pad3, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , __A21_1__C45M, __A21_1__C46M, __A21_1__C57A, __A21_1__C60A, net_U21015_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21016(net_U21016_Pad1, __A21_1__30SUM, __A21_1__50SUM, CAD1, __A21_1__RSCT_n, net_R21001_Pad2, GND, __A21_1__RSCT_n, net_R21002_Pad2, CAD2, __A21_1__RSCT_n, net_R21003_Pad2, CAD3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21017(CAD4, __A21_1__RSCT_n, net_U21016_Pad1, CAD5, __A21_1__RSCT_n, net_R21006_Pad2, GND, __A21_1__RSCT_n, net_R21007_Pad2, CAD6, __A21_1__C45P, __A21_1__C46P, net_U21017_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21018(C31A, __A21_1__C47A, C51A, C52A, C53A, net_U21014_Pad11, GND, net_U21014_Pad13, C54A, C55A, __A21_1__C56A, net_U21014_Pad9, C50A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U21019(net_U21019_Pad1, INCSET_n, net_U21015_Pad13, net_U21019_Pad4, INCSET_n, net_U21017_Pad13, GND, INCSET_n, net_R21008_Pad2, net_U21019_Pad10, net_U21019_Pad1, __A21_1__SHINC, SHINC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21020(__A21_1__SHINC, SHINC_n, T12A, SHANC_n, net_U21019_Pad4, __A21_1__SHANC, GND, SHANC_n, T12A, __A21_1__SHANC, net_U21019_Pad10, DINC, __A21_1__DINCNC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21021(DINC, __A21_1__DINCNC_n, T12A, net_U21021_Pad4, INCSET_n, net_R21009_Pad2, GND, net_U21021_Pad4, PINC, __A21_1__PINC_n, __A21_1__PINC_n, T12, PINC, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21022(net_U21022_Pad1, C24A, C25A, C26A, C27A,  , GND,  , C30A, C37P, C40P, C41P, net_U21022_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21023(net_U21022_Pad1, net_R21009_Pad2, net_U21022_Pad13, net_R21009_Pad2, net_U21023_Pad5, net_R21009_Pad2, GND, net_R21010_Pad2, net_U21023_Pad9, net_R21010_Pad2, net_U21023_Pad11, net_R21011_Pad2, net_U21023_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U21024(__A21_1__C42P, __A21_1__C43P, __A21_1__C42M, __A21_1__C43M, __A21_1__C44M, net_U21023_Pad9, GND, net_U21023_Pad11, C37M, C40M, C41M, net_U21023_Pad5, __A21_1__C44P, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21025(net_U21025_Pad1, INCSET_n, net_R21010_Pad2, __A21_1__MINC_n, net_U21025_Pad1, MINC, GND, __A21_1__MINC_n, T12A, MINC, C35P, C36P, net_U21025_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21026(C32P, C33P, C32M, C33M, C34M, net_U21026_Pad6, GND,  ,  ,  ,  , net_U21023_Pad13, C34P, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21027(net_U21025_Pad13, net_R21011_Pad2, net_U21026_Pad6, net_R21012_Pad2, net_U21027_Pad5, net_R21012_Pad2, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21028(net_U21028_Pad1, INCSET_n, net_R21011_Pad2, __A21_1__PCDU_n, net_U21028_Pad1, PCDU, GND, __A21_1__PCDU_n, T12A, PCDU, C35M, C36M, net_U21027_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21029(net_U21029_Pad1, INCSET_n, net_R21012_Pad2, __A21_1__MCDU_n, net_U21029_Pad1, MCDU, GND, __A21_1__MCDU_n, T12A, MCDU, net_U21029_Pad11, __A21_3__C43R, net_U21029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21030(net_U21030_Pad1, BMAGXP, net_U21030_Pad3, net_U21030_Pad3, net_U21030_Pad1, __A21_3__C42R, GND, BMAGXM, net_U21030_Pad13, net_U21030_Pad10, net_U21030_Pad10, __A21_3__C42R, net_U21030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U21031(BKTF_n, net_U21031_Pad2, RSSB, net_U21031_Pad4, net_U21031_Pad5, __A21_3__CG15, GND, CTROR, CTROR_n, net_U21031_Pad10, RSSB, net_U21031_Pad12, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21032(net_U21032_Pad1, net_U21030_Pad3, net_U21030_Pad13, net_U21032_Pad4, net_U21031_Pad2, net_U21032_Pad1, GND, net_U21032_Pad4, net_U21032_Pad13, net_U21032_Pad10, net_U21032_Pad10, __A21_3__C42R, net_U21032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21033(__A21_1__C42A, CG13, net_U21032_Pad10, net_U21029_Pad11, BMAGYP, net_U21029_Pad13, GND, __A21_1__SHINC, __A21_1__SHANC, SHIFT_n, BMAGYM, net_U21033_Pad12, net_U21033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21034(net_U21031_Pad4, CA4_n, net_U21030_Pad1, CA4_n, CXB2_n, __A21_1__C42P, GND, __A21_1__C42M, net_U21030_Pad10, CA4_n, CXB2_n, __A21_3__C42R, CXB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21035(net_U21033_Pad12, net_U21033_Pad13, __A21_3__C43R, net_U21035_Pad4, net_U21029_Pad13, net_U21033_Pad12, GND, net_U21031_Pad2, net_U21035_Pad4, net_U21035_Pad10, net_U21035_Pad10, net_U21035_Pad12, net_U21035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21036(net_U21035_Pad12, net_U21035_Pad13, __A21_3__C43R, net_U21036_Pad12, EMSD, net_U21036_Pad10, GND, net_U21036_Pad12, __A21_3__C56R, net_U21036_Pad10, net_U21031_Pad2, net_U21036_Pad12, net_U21036_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21037(net_U21031_Pad4, CA4_n, net_U21029_Pad11, CA4_n, CXB3_n, __A21_1__C43P, GND, __A21_1__C43M, net_U21033_Pad13, CA4_n, CXB3_n, __A21_3__C43R, CXB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21038(CG13, net_U21032_Pad13, CG13, net_U21032_Pad13, net_U21035_Pad12, net_U21031_Pad5, GND, __A21_3__C56R, net_U21031_Pad4, CA5_n, CXB6_n, __A21_1__C43A, net_U21035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21039(net_U21039_Pad1, net_U21036_Pad13, net_U21039_Pad3, net_U21039_Pad3, net_U21039_Pad1, __A21_3__C56R, GND, CG23, net_U21039_Pad1, __A21_1__C56A, OTLNKM, net_U21039_Pad12, net_U21039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21040(net_U21039_Pad12, net_U21039_Pad13, __A21_3__C57R, net_U21040_Pad4, net_U21031_Pad2, net_U21039_Pad13, GND, net_U21040_Pad4, net_U21040_Pad13, net_U21040_Pad10, net_U21040_Pad10, __A21_3__C57R, net_U21040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21041(net_U21031_Pad4, CA5_n, CG23, net_U21039_Pad3, net_U21040_Pad10, __A21_1__C57A, GND, __A21_3__C60R, net_U21031_Pad4, CA6_n, CXB0_n, __A21_3__C57R, CXB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U21042(net_U21042_Pad1, ALTM, net_U21042_Pad3, net_U21042_Pad3, net_U21042_Pad1, __A21_3__C60R, GND, net_U21031_Pad2, net_U21042_Pad1, net_U21042_Pad10, net_U21042_Pad10, net_U21042_Pad12, net_U21042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21043(net_U21042_Pad12, net_U21042_Pad13, __A21_3__C60R, net_U21043_Pad4, BMAGZP, net_U21043_Pad10, GND, net_U21043_Pad4, __A21_3__C44R, net_U21043_Pad10, BMAGZM, net_U21043_Pad12, net_U21043_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21044(__A21_1__C60A, CG23, net_U21039_Pad3, net_U21040_Pad13, net_U21042_Pad13,  , GND,  , CG23, net_U21039_Pad3, net_U21040_Pad13, net_U21042_Pad12, CTROR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21045(net_U21043_Pad12, net_U21043_Pad13, __A21_3__C44R, net_U21045_Pad4, net_U21043_Pad10, net_U21043_Pad12, net_U21045_Pad7, net_U21031_Pad12, net_U21045_Pad4, net_U21045_Pad10, net_U21045_Pad10, net_U21045_Pad12, net_U21045_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21046(net_U21045_Pad12, net_U21045_Pad13, __A21_3__C44R, __A21_1__C44A, __A21_3__CG15, net_U21045_Pad13, GND, INLNKP, net_U21046_Pad13, net_U21046_Pad10, net_U21046_Pad10, C45R, net_U21046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21047(net_U21031_Pad10, CA4_n, net_U21043_Pad4, CA4_n, CXB4_n, __A21_1__C44P, GND, __A21_1__C44M, net_U21043_Pad13, CA4_n, CXB4_n, __A21_3__C44R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21048(net_U21048_Pad1, INLNKM, net_U21048_Pad3, net_U21048_Pad3, net_U21048_Pad1, C45R, GND, net_U21046_Pad13, net_U21048_Pad3, net_U21048_Pad10, net_U21031_Pad12, net_U21048_Pad10, net_U21048_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21049(net_U21049_Pad1, net_U21048_Pad13, net_U21049_Pad3, net_U21049_Pad3, net_U21049_Pad1, C45R, GND, RNRADP, net_U21049_Pad13, net_U21049_Pad10, net_U21049_Pad10, __A21_3__C46R, net_U21049_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21050(net_U21031_Pad10, CA4_n, net_U21046_Pad10, CA4_n, CXB5_n, __A21_1__C45P, GND, __A21_1__C45M, net_U21048_Pad1, CA4_n, CXB5_n, C45R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21051(__A21_3__CG15, net_U21045_Pad12, __A21_3__CG15, net_U21045_Pad12, net_U21049_Pad3, net_U21051_Pad6, GND, __A21_3__C46R, net_U21031_Pad10, CA4_n, CXB6_n, __A21_1__C45A, net_U21049_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21052(net_U21051_Pad6, __A21_3__CG16, net_U21052_Pad3, CG26, XB3, CXB3_n, GND, CXB4_n, XB4, CXB5_n, XB5, CXB6_n, XB6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21053(net_U21053_Pad1, net_U21031_Pad12, net_U21053_Pad3, net_U21053_Pad12, net_U21053_Pad1, net_U21053_Pad10, GND, net_U21053_Pad12, __A21_3__C46R, net_U21053_Pad10, __A21_3__CG16, net_U21053_Pad12, __A21_1__C46A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21054(net_U21054_Pad1, RNRADM, net_U21054_Pad3, net_U21054_Pad3, net_U21054_Pad1, __A21_3__C46R, GND, net_U21049_Pad13, net_U21054_Pad3, net_U21053_Pad3, net_U21054_Pad11, net_U21054_Pad12, net_U21054_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21055(net_U21054_Pad12, net_U21054_Pad13, __A21_3__C47R, net_U21055_Pad12, GYROD, net_U21055_Pad10, GND, net_U21055_Pad12, __A21_3__C47R, net_U21055_Pad10, net_U21031_Pad12, net_U21055_Pad12, net_U21054_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21056(net_U21049_Pad10, CA4_n, CA4_n, CXB6_n, net_U21054_Pad1, __A21_1__C46M, GND, __A21_3__C47R, net_U21031_Pad10, CA4_n, CXB7_n, __A21_1__C46P, CXB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21057(__A21_3__CG16, net_U21053_Pad10, __A21_3__CG16, net_U21053_Pad10, net_U21054_Pad12, net_U21052_Pad3, GND,  ,  ,  ,  , __A21_1__C47A, net_U21054_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21058(XB7, CXB7_n, OCTAD2, CA2_n, OCTAD3, CA3_n, GND, CA4_n, OCTAD4, CA5_n, OCTAD5, CA6_n, OCTAD6, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21059(SHIFT_n, SHIFT, RSCT, __A21_1__RSCT_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule