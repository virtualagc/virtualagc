`timescale 1ns/1ps
`default_nettype none

module counter_cell_ii(SIM_RST, SIM_CLK, p4VSW, GND, T12, T12A, INCSET_n, RSCT, BKTF_n, RSSB, BMAGXP, BMAGXM, BMAGYP, BMAGYM, EMSD, OTLNKM, ALTM, BMAGZP, BMAGZM, INLNKP, INLNKM, RNRADP, RNRADM, GYROD, XB0, XB1, XB2, XB3, XB4, XB5, XB6, XB7, OCTAD2, OCTAD3, OCTAD4, OCTAD5, OCTAD6, CG13, CG23, C24A, C25A, C26A, C27A, C30A, C31A, C32A, C32P, C32M, C33A, C33P, C33M, C34A, C34P, C34M, C35A, C35P, C35M, C36A, C36P, C36M, C37A, C37P, C37M, C40A, C40P, C40M, C41A, C41P, C41M, C50A, C51A, C52A, C53A, C54A, C55A, CA2_n, CA3_n, CA4_n, CA5_n, CA6_n, CXB0_n, CXB1_n, CXB2_n, CXB3_n, CXB4_n, CXB5_n, CXB6_n, CXB7_n, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CG26, C45R, PINC, MINC, DINC, DINC_n, PCDU, MCDU, SHINC_n, SHANC_n, SHIFT, SHIFT_n, CTROR, CTROR_n);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire ALTM;
    input wire BKTF_n;
    input wire BMAGXM;
    input wire BMAGXP;
    input wire BMAGYM;
    input wire BMAGYP;
    input wire BMAGZM;
    input wire BMAGZP;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C31A;
    input wire C32A;
    input wire C32M;
    input wire C32P;
    input wire C33A;
    input wire C33M;
    input wire C33P;
    input wire C34A;
    input wire C34M;
    input wire C34P;
    input wire C35A;
    input wire C35M;
    input wire C35P;
    input wire C36A;
    input wire C36M;
    input wire C36P;
    input wire C37A;
    input wire C37M;
    input wire C37P;
    input wire C40A;
    input wire C40M;
    input wire C40P;
    input wire C41A;
    input wire C41M;
    input wire C41P;
    output wire C45R;
    input wire C50A;
    input wire C51A;
    input wire C52A;
    input wire C53A;
    input wire C54A;
    input wire C55A;
    output wire CA2_n;
    output wire CA3_n;
    output wire CA4_n;
    output wire CA5_n;
    output wire CA6_n;
    output wire CAD1;
    output wire CAD2;
    output wire CAD3;
    output wire CAD4;
    output wire CAD5;
    output wire CAD6;
    input wire CG13;
    input wire CG23;
    output wire CG26;
    output wire CTROR;
    output wire CTROR_n;
    output wire CXB0_n;
    output wire CXB1_n;
    output wire CXB2_n;
    output wire CXB3_n;
    output wire CXB4_n;
    output wire CXB5_n;
    output wire CXB6_n;
    output wire CXB7_n;
    output wire DINC;
    output wire DINC_n;
    input wire EMSD;
    input wire GYROD;
    input wire INCSET_n;
    input wire INLNKM;
    input wire INLNKP;
    output wire MCDU;
    output wire MINC;
    input wire OCTAD2;
    input wire OCTAD3;
    input wire OCTAD4;
    input wire OCTAD5;
    input wire OCTAD6;
    input wire OTLNKM;
    output wire PCDU;
    output wire PINC;
    input wire RNRADM;
    input wire RNRADP;
    input wire RSCT;
    input wire RSSB;
    output wire SHANC_n;
    output wire SHIFT;
    output wire SHIFT_n;
    output wire SHINC_n;
    input wire T12;
    input wire T12A;
    input wire XB0;
    input wire XB1;
    input wire XB2;
    input wire XB3;
    input wire XB4;
    input wire XB5;
    input wire XB6;
    input wire XB7;
    wire __A21_1__30SUM;
    wire __A21_1__32004K; //FPGA#wand
    wire __A21_1__50SUM;
    wire __A21_1__C42A;
    wire __A21_1__C42M;
    wire __A21_1__C42P;
    wire __A21_1__C43A;
    wire __A21_1__C43M;
    wire __A21_1__C43P;
    wire __A21_1__C44A;
    wire __A21_1__C44M;
    wire __A21_1__C44P;
    wire __A21_1__C45A;
    wire __A21_1__C45M;
    wire __A21_1__C45P;
    wire __A21_1__C46A;
    wire __A21_1__C46M;
    wire __A21_1__C46P;
    wire __A21_1__C47A;
    wire __A21_1__C56A;
    wire __A21_1__C57A;
    wire __A21_1__C60A;
    wire __A21_1__DINCNC_n;
    wire __A21_1__MCDU_n;
    wire __A21_1__MINC_n;
    wire __A21_1__PCDU_n;
    wire __A21_1__PINC_n;
    wire __A21_1__RSCT_n;
    wire __A21_1__SHANC;
    wire __A21_1__SHINC;
    wire __A21_3__C42R;
    wire __A21_3__C43R;
    wire __A21_3__C44R;
    wire __A21_3__C46R;
    wire __A21_3__C47R;
    wire __A21_3__C56R;
    wire __A21_3__C57R;
    wire __A21_3__C60R;
    wire __A21_3__CG15;
    wire __A21_3__CG16;
    wire __A21_NET_133;
    wire __A21_NET_134;
    wire __A21_NET_136;
    wire __A21_NET_140;
    wire __A21_NET_141; //FPGA#wand
    wire __A21_NET_142;
    wire __A21_NET_143;
    wire __A21_NET_144;
    wire __A21_NET_145; //FPGA#wand
    wire __A21_NET_146; //FPGA#wand
    wire __A21_NET_147; //FPGA#wand
    wire __A21_NET_148;
    wire __A21_NET_149;
    wire __A21_NET_151;
    wire __A21_NET_152; //FPGA#wand
    wire __A21_NET_153; //FPGA#wand
    wire __A21_NET_154;
    wire __A21_NET_156;
    wire __A21_NET_157;
    wire __A21_NET_159; //FPGA#wand
    wire __A21_NET_160;
    wire __A21_NET_161;
    wire __A21_NET_162; //FPGA#wand
    wire __A21_NET_163;
    wire __A21_NET_164;
    wire __A21_NET_165;
    wire __A21_NET_166;
    wire __A21_NET_168;
    wire __A21_NET_172;
    wire __A21_NET_173; //FPGA#wand
    wire __A21_NET_174;
    wire __A21_NET_178;
    wire __A21_NET_179;
    wire __A21_NET_184;
    wire __A21_NET_185;
    wire __A21_NET_187; //FPGA#wand
    wire __A21_NET_188;
    wire __A21_NET_193;
    wire __A21_NET_194;
    wire __A21_NET_199;
    wire __A21_NET_200;
    wire __A21_NET_203;
    wire __A21_NET_204;
    wire __A21_NET_205;
    wire __A21_NET_212;
    wire __A21_NET_215;
    wire __A21_NET_216;
    wire __A21_NET_219;
    wire __A21_NET_224;
    wire __A21_NET_225;
    wire __A21_NET_226;
    wire __A21_NET_227;
    wire __A21_NET_228;
    wire __A21_NET_229; //FPGA#wand
    wire __A21_NET_232;
    wire __A21_NET_233;
    wire __A21_NET_234;
    wire __A21_NET_235;
    wire __A21_NET_236;
    wire __A21_NET_237;
    wire __A21_NET_238;
    wire __A21_NET_239;
    wire __A21_NET_240;
    wire __A21_NET_241;
    wire __A21_NET_242;
    wire __A21_NET_243;
    wire __A21_NET_244;
    wire __A21_NET_245;
    wire __A21_NET_246;
    wire __A21_NET_247;
    wire __A21_NET_248;
    wire __A21_NET_249;
    wire __A21_NET_250;
    wire __A21_NET_251;
    wire __A21_NET_252;
    wire __A21_NET_253;
    wire __A21_NET_254;
    wire __A21_NET_255;
    wire __A21_NET_256;
    wire __A21_NET_257;
    wire __A21_NET_258;
    wire __A21_NET_259;
    wire __A21_NET_260;
    wire __A21_NET_261;
    wire __A21_NET_262;
    wire __A21_NET_263;
    wire __A21_NET_264;
    wire __A21_NET_265;
    wire __A21_NET_266;
    wire __A21_NET_267;
    wire __A21_NET_268;
    wire __A21_NET_269;
    wire __A21_NET_271;
    wire __A21_NET_272;
    wire __A21_NET_273;
    wire __A21_NET_274;
    wire __A21_NET_275;
    wire __A21_NET_276;
    wire __A21_NET_277;
    wire __A21_NET_278;
    wire __A21_NET_279;
    wire __A21_NET_280;
    wire __A21_NET_281;
    wire __A21_NET_282;
    wire __A21_NET_283;
    wire __A21_NET_284;
    wire __A21_NET_285;
    wire __A21_NET_286;
    wire __A21_NET_287;
    wire __A21_NET_288;
    wire __A21_NET_289;
    wire __A21_NET_290;
    wire __A21_NET_292;
    wire __A21_NET_300;
    wire __A21_NET_301;
    wire __A21_NET_302;
    wire __A21_NET_304;
    wire __A21_NET_305;
    wire __A21_NET_306;
    wire __A21_NET_307;
    wire __A21_NET_308;
    wire __A21_NET_71;

    pullup R21001(__A21_NET_152);
    pullup R21002(__A21_NET_153);
    pullup R21003(__A21_NET_147);
    pullup R21004(__A21_1__32004K);
    pullup R21005(__A21_NET_173);
    pullup R21006(__A21_NET_146);
    pullup R21007(__A21_NET_187);
    pullup R21008(__A21_NET_229);
    pullup R21009(__A21_NET_141);
    pullup R21010(__A21_NET_145);
    pullup R21011(__A21_NET_159);
    pullup R21012(__A21_NET_162);
    U74HC4002 U21001(__A21_NET_205, C25A, C27A, C31A, C33A,  , GND,  , C35A, C37A, C41A, __A21_1__C43A, __A21_NET_204, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21002(__A21_NET_205, __A21_NET_152, __A21_NET_204, __A21_NET_152, __A21_NET_199, __A21_NET_152, GND, __A21_NET_152, __A21_NET_200, __A21_NET_153, __A21_NET_203, __A21_NET_153, __A21_NET_219, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21003(__A21_NET_199, __A21_1__C45A, __A21_1__C47A, C51A, C53A,  , GND,  , C26A, C27A, C32A, C33A, __A21_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21004(__A21_NET_200, C55A, __A21_1__C57A, __A21_NET_225, __A21_1__C56A, __A21_1__C57A, GND, __A21_1__30SUM, __A21_1__C60A, __A21_NET_188, __A21_1__50SUM, __A21_1__C60A, __A21_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21005(__A21_NET_219, C36A, C37A, __A21_1__C42A, __A21_1__C43A,  , GND,  , __A21_1__C46A, __A21_1__C47A, C52A, C53A, __A21_NET_224, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21006(__A21_NET_224, __A21_NET_153, __A21_NET_225, __A21_NET_153, __A21_NET_212, __A21_NET_147, GND, __A21_NET_147, __A21_NET_215, __A21_NET_147, __A21_NET_216, __A21_NET_147, __A21_NET_178, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21007(__A21_NET_212, C24A, C25A, C26A, C27A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21008(__A21_NET_216, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_178, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21009(__A21_NET_179, C30A, C31A, C32A, C33A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21010(__A21_NET_179, __A21_1__32004K, __A21_NET_184, __A21_1__32004K, __A21_NET_168, __A21_NET_173, GND, __A21_NET_173, __A21_NET_172, __A21_NET_146, __A21_NET_174, __A21_NET_146, __A21_NET_188, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC04 U21011(__A21_1__32004K, __A21_1__30SUM, __A21_NET_173, __A21_1__50SUM, DINC, DINC_n, GND, CXB0_n, XB0, CXB1_n, XB1, CXB2_n, XB2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21012(__A21_NET_168, C50A, C51A, C52A, C53A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_172, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21013(__A21_NET_174, C24A, C25A, C26A, C27A,  , GND,  , C40A, C41A, __A21_1__C42A, __A21_1__C43A, __A21_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21014(__A21_NET_193, __A21_NET_187, __A21_NET_194, __A21_NET_187, __A21_NET_185, __A21_NET_187, GND, __A21_NET_229, __A21_NET_228, __A21_NET_229, __A21_NET_227, __A21_NET_229, __A21_NET_226, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21015(__A21_NET_194, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , __A21_1__C45M, __A21_1__C46M, __A21_1__C57A, __A21_1__C60A, __A21_NET_148, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21016(__A21_NET_151, __A21_1__30SUM, __A21_1__50SUM, CAD1, __A21_1__RSCT_n, __A21_NET_152, GND, __A21_1__RSCT_n, __A21_NET_153, CAD2, __A21_1__RSCT_n, __A21_NET_147, CAD3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21017(CAD4, __A21_1__RSCT_n, __A21_NET_151, CAD5, __A21_1__RSCT_n, __A21_NET_146, GND, __A21_1__RSCT_n, __A21_NET_187, CAD6, __A21_1__C45P, __A21_1__C46P, __A21_NET_149, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21018(C31A, __A21_1__C47A, C51A, C52A, C53A, __A21_NET_227, GND, __A21_NET_226, C54A, C55A, __A21_1__C56A, __A21_NET_228, C50A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U21019(__A21_NET_156, INCSET_n, __A21_NET_148, __A21_NET_157, INCSET_n, __A21_NET_149, GND, INCSET_n, __A21_NET_229, __A21_NET_154, __A21_NET_156, __A21_1__SHINC, SHINC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21020(__A21_1__SHINC, SHINC_n, T12A, SHANC_n, __A21_NET_157, __A21_1__SHANC, GND, SHANC_n, T12A, __A21_1__SHANC, __A21_NET_154, DINC, __A21_1__DINCNC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21021(DINC, __A21_1__DINCNC_n, T12A, __A21_NET_133, INCSET_n, __A21_NET_141, GND, __A21_NET_133, PINC, __A21_1__PINC_n, __A21_1__PINC_n, T12, PINC, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21022(__A21_NET_136, C24A, C25A, C26A, C27A,  , GND,  , C30A, C37P, C40P, C41P, __A21_NET_140, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21023(__A21_NET_136, __A21_NET_141, __A21_NET_140, __A21_NET_141, __A21_NET_134, __A21_NET_141, GND, __A21_NET_145, __A21_NET_144, __A21_NET_145, __A21_NET_142, __A21_NET_159, __A21_NET_164, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U21024(__A21_1__C42P, __A21_1__C43P, __A21_1__C42M, __A21_1__C43M, __A21_1__C44M, __A21_NET_144, GND, __A21_NET_142, C37M, C40M, C41M, __A21_NET_134, __A21_1__C44P, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21025(__A21_NET_143, INCSET_n, __A21_NET_145, __A21_1__MINC_n, __A21_NET_143, MINC, GND, __A21_1__MINC_n, T12A, MINC, C35P, C36P, __A21_NET_160, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21026(C32P, C33P, C32M, C33M, C34M, __A21_NET_161, GND,  ,  ,  ,  , __A21_NET_164, C34P, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21027(__A21_NET_160, __A21_NET_159, __A21_NET_161, __A21_NET_162, __A21_NET_163, __A21_NET_162, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21028(__A21_NET_166, INCSET_n, __A21_NET_159, __A21_1__PCDU_n, __A21_NET_166, PCDU, GND, __A21_1__PCDU_n, T12A, PCDU, C35M, C36M, __A21_NET_163, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21029(__A21_NET_165, INCSET_n, __A21_NET_162, __A21_1__MCDU_n, __A21_NET_165, MCDU, GND, __A21_1__MCDU_n, T12A, MCDU, __A21_NET_249, __A21_3__C43R, __A21_NET_252, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21030(__A21_NET_300, BMAGXP, __A21_NET_305, __A21_NET_305, __A21_NET_300, __A21_3__C42R, GND, BMAGXM, __A21_NET_304, __A21_NET_302, __A21_NET_302, __A21_3__C42R, __A21_NET_304, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U21031(BKTF_n, __A21_NET_301, RSSB, __A21_NET_276, __A21_NET_262, __A21_3__CG15, GND, CTROR, CTROR_n, __A21_NET_244, RSSB, __A21_NET_241, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21032(__A21_NET_306, __A21_NET_305, __A21_NET_304, __A21_NET_307, __A21_NET_301, __A21_NET_306, GND, __A21_NET_307, __A21_NET_261, __A21_NET_308, __A21_NET_308, __A21_3__C42R, __A21_NET_261, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21033(__A21_1__C42A, CG13, __A21_NET_308, __A21_NET_249, BMAGYP, __A21_NET_252, GND, __A21_1__SHINC, __A21_1__SHANC, SHIFT_n, BMAGYM, __A21_NET_253, __A21_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21034(__A21_NET_276, CA4_n, __A21_NET_300, CA4_n, CXB2_n, __A21_1__C42P, GND, __A21_1__C42M, __A21_NET_302, CA4_n, CXB2_n, __A21_3__C42R, CXB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21035(__A21_NET_253, __A21_NET_250, __A21_3__C43R, __A21_NET_254, __A21_NET_252, __A21_NET_253, GND, __A21_NET_301, __A21_NET_254, __A21_NET_256, __A21_NET_256, __A21_NET_255, __A21_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21036(__A21_NET_255, __A21_NET_251, __A21_3__C43R, __A21_NET_264, EMSD, __A21_NET_263, GND, __A21_NET_264, __A21_3__C56R, __A21_NET_263, __A21_NET_301, __A21_NET_264, __A21_NET_258, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21037(__A21_NET_276, CA4_n, __A21_NET_249, CA4_n, CXB3_n, __A21_1__C43P, GND, __A21_1__C43M, __A21_NET_250, CA4_n, CXB3_n, __A21_3__C43R, CXB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21038(CG13, __A21_NET_261, CG13, __A21_NET_261, __A21_NET_255, __A21_NET_262, GND, __A21_3__C56R, __A21_NET_276, CA5_n, CXB6_n, __A21_1__C43A, __A21_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21039(__A21_NET_257, __A21_NET_258, __A21_NET_236, __A21_NET_236, __A21_NET_257, __A21_3__C56R, GND, CG23, __A21_NET_257, __A21_1__C56A, OTLNKM, __A21_NET_259, __A21_NET_260, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21040(__A21_NET_259, __A21_NET_260, __A21_3__C57R, __A21_NET_238, __A21_NET_301, __A21_NET_260, GND, __A21_NET_238, __A21_NET_245, __A21_NET_237, __A21_NET_237, __A21_3__C57R, __A21_NET_245, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21041(__A21_NET_276, CA5_n, CG23, __A21_NET_236, __A21_NET_237, __A21_1__C57A, GND, __A21_3__C60R, __A21_NET_276, CA6_n, CXB0_n, __A21_3__C57R, CXB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U21042(__A21_NET_234, ALTM, __A21_NET_239, __A21_NET_239, __A21_NET_234, __A21_3__C60R, GND, __A21_NET_301, __A21_NET_234, __A21_NET_235, __A21_NET_235, __A21_NET_233, __A21_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21043(__A21_NET_233, __A21_NET_232, __A21_3__C60R, __A21_NET_288, BMAGZP, __A21_NET_246, GND, __A21_NET_288, __A21_3__C44R, __A21_NET_246, BMAGZM, __A21_NET_247, __A21_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21044(__A21_1__C60A, CG23, __A21_NET_236, __A21_NET_245, __A21_NET_232,  , GND,  , CG23, __A21_NET_236, __A21_NET_245, __A21_NET_233, CTROR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21045(__A21_NET_247, __A21_NET_248, __A21_3__C44R, __A21_NET_240, __A21_NET_246, __A21_NET_247, __A21_NET_71, __A21_NET_241, __A21_NET_240, __A21_NET_243, __A21_NET_243, __A21_NET_292, __A21_NET_242, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21046(__A21_NET_292, __A21_NET_242, __A21_3__C44R, __A21_1__C44A, __A21_3__CG15, __A21_NET_242, GND, INLNKP, __A21_NET_283, __A21_NET_289, __A21_NET_289, C45R, __A21_NET_283, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21047(__A21_NET_244, CA4_n, __A21_NET_288, CA4_n, CXB4_n, __A21_1__C44P, GND, __A21_1__C44M, __A21_NET_248, CA4_n, CXB4_n, __A21_3__C44R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21048(__A21_NET_282, INLNKM, __A21_NET_281, __A21_NET_281, __A21_NET_282, C45R, GND, __A21_NET_283, __A21_NET_281, __A21_NET_284, __A21_NET_241, __A21_NET_284, __A21_NET_287, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21049(__A21_NET_286, __A21_NET_287, __A21_NET_285, __A21_NET_285, __A21_NET_286, C45R, GND, RNRADP, __A21_NET_290, __A21_NET_275, __A21_NET_275, __A21_3__C46R, __A21_NET_290, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21050(__A21_NET_244, CA4_n, __A21_NET_289, CA4_n, CXB5_n, __A21_1__C45P, GND, __A21_1__C45M, __A21_NET_282, CA4_n, CXB5_n, C45R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21051(__A21_3__CG15, __A21_NET_292, __A21_3__CG15, __A21_NET_292, __A21_NET_285, __A21_NET_277, GND, __A21_3__C46R, __A21_NET_244, CA4_n, CXB6_n, __A21_1__C45A, __A21_NET_286, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21052(__A21_NET_277, __A21_3__CG16, __A21_NET_278, CG26, XB3, CXB3_n, GND, CXB4_n, XB4, CXB5_n, XB5, CXB6_n, XB6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21053(__A21_NET_273, __A21_NET_241, __A21_NET_280, __A21_NET_272, __A21_NET_273, __A21_NET_271, GND, __A21_NET_272, __A21_3__C46R, __A21_NET_271, __A21_3__CG16, __A21_NET_272, __A21_1__C46A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21054(__A21_NET_274, RNRADM, __A21_NET_279, __A21_NET_279, __A21_NET_274, __A21_3__C46R, GND, __A21_NET_290, __A21_NET_279, __A21_NET_280, __A21_NET_269, __A21_NET_265, __A21_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21055(__A21_NET_265, __A21_NET_268, __A21_3__C47R, __A21_NET_267, GYROD, __A21_NET_266, GND, __A21_NET_267, __A21_3__C47R, __A21_NET_266, __A21_NET_241, __A21_NET_267, __A21_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21056(__A21_NET_275, CA4_n, CA4_n, CXB6_n, __A21_NET_274, __A21_1__C46M, GND, __A21_3__C47R, __A21_NET_244, CA4_n, CXB7_n, __A21_1__C46P, CXB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21057(__A21_3__CG16, __A21_NET_271, __A21_3__CG16, __A21_NET_271, __A21_NET_265, __A21_NET_278, GND,  ,  ,  ,  , __A21_1__C47A, __A21_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21058(XB7, CXB7_n, OCTAD2, CA2_n, OCTAD3, CA3_n, GND, CA4_n, OCTAD4, CA5_n, OCTAD5, CA6_n, OCTAD6, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21059(SHIFT_n, SHIFT, RSCT, __A21_1__RSCT_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule