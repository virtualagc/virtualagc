// Verilog testbench created by dumbTestbench.py
`timescale 1ns / 1ps

module agc;

parameter GATE_DELAY = 20;
`include "tb-2003200.v"

reg BLKUPL_ = 1, BMGXM = 0, BMGXP = 0, BMGYM = 0, BMGYP = 0, BMGZM = 0,
  BMGZP = 0, CAURST = 0, CDUFAL = 0, CDUXM = 0, CDUXP = 0, CDUYM = 0, CDUYP = 0,
  CDUZM = 0, CDUZP = 0, CGA1 = 0, CGA10 = 0, CGA11 = 0, CGA12 = 0, CGA13 = 0,
  CGA14 = 0, CGA15 = 0, CGA16 = 0, CGA17 = 0, CGA18 = 0, CGA19 = 0, CGA2 = 0,
  CGA20 = 0, CGA21 = 0, CGA22 = 0, CGA23 = 0, CGA24 = 0, CGA3 = 0, CGA4 = 0,
  CGA5 = 0, CGA6 = 0, CGA7 = 0, CGA8 = 0, CGA9 = 0, CTLSAT = 0, FLTOUT = 0,
  FREFUN = 0, GATEX_ = 1, GATEY_ = 1, GATEZ_ = 1, GCAPCL = 0, GUIREL = 0,
  HOLFUN = 0, IMUCAG = 0, IMUFAL = 0, IMUOPR = 0, IN3008 = 0, IN3212 = 0,
  IN3213 = 0, IN3214 = 0, IN3216 = 0, IN3301 = 0, ISSTOR = 0, LEMATT = 0,
  LFTOFF = 0, LRIN0 = 0, LRIN1 = 0, LRRLSC = 0, LVDAGD = 0, MAINRS = 0,
  MANRmP = 0, MANRmR = 0, MANRmY = 0, MANRpP = 0, MANRpR = 0, MANRpY = 0,
  MARK = 0, MKEY1 = 0, MKEY2 = 0, MKEY3 = 0, MKEY4 = 0, MKEY5 = 0, MNIMmP = 0,
  MNIMmR = 0, MNIMmY = 0, MNIMpP = 0, MNIMpR = 0, MNIMpY = 0, MRKREJ = 0,
  MRKRST = 0, NAVRST = 0, NHVFAL = 0, NKEY1 = 0, NKEY2 = 0, NKEY3 = 0,
  NKEY4 = 0, NKEY5 = 0, OPCDFL = 0, OPMSW2 = 0, OPMSW3 = 0, PCHGOF = 0,
  ROLGOF = 0, RRIN0 = 0, RRIN1 = 0, RRPONA = 0, RRRLSC = 0, S4BSAB = 0,
  SBYBUT = 0, SCAFAL = 0, SHAFTM = 0, SHAFTP = 0, SIGNX = 0, SIGNY = 0,
  SIGNZ = 0, SMSEPR = 0, SPSRDY = 0, STRPRS = 0, STRT2 = 0, TEMPIN = 0,
  TRANmX = 0, TRANmY = 0, TRANmZ = 0, TRANpX = 0, TRANpY = 0, TRANpZ = 0,
  TRNM = 0, TRNP = 0, TRST10 = 0, TRST9 = 0, ULLTHR = 0, UPL0 = 0, UPL1 = 0,
  VFAIL = 0, XLNK0 = 0, XLNK1 = 0, ZEROP = 0, d2FSFAL = 0, p4SW = 0;

wire A01_, A02_, A03_, A04_, A05_, A06_, A07_, A08_, A09_, A10_, A11_,
  A12_, A13_, A14_, A15_, A16_, A2XG_, A2X_, AD0, ADS0, ADVCTR, AGCWAR,
  ALGA, ALRT0, ALRT1, ALT0, ALT1, ALTEST, ALTM, ALTSNC, AUG0, AUG0_, B15X,
  BBK1, BBK2, BBK3, BK16, BKTF_, BLKUPL, BMAGXM, BMAGXP, BMAGYM, BMAGYP,
  BMAGZM, BMAGZP, BMF0, BMF0_, BOTHX, BOTHY, BOTHZ, BR1, BR12B, BR12B_,
  BR1B2, BR1B2B, BR1B2B_, BR1B2_, BR1_, BR2, BR2_, BRDIF_, BRXP3, BSYNC_,
  BXVX, BZF0, BZF0_, C24A, C24R, C25A, C25R, C26A, C26R, C27A, C27R, C30A,
  C30R, C31A, C31R, C32A, C32M, C32P, C32R, C33A, C33M, C33P, C33R, C34A,
  C34M, C34P, C34R, C35A, C35M, C35P, C35R, C36A, C36M, C36P, C36R, C37A,
  C37M, C37P, C37R, C40A, C40M, C40P, C40R, C41A, C41M, C41P, C41R, C42A,
  C42M, C42P, C42R, C43A, C43M, C43P, C43R, C44A, C44M, C44P, C44R, C45A,
  C45M, C45P, C45R, C45R_, C46A, C46M, C46P, C46R, C47A, C47R, C50A, C50R,
  C51A, C51R, C52A, C52R, C53A, C53R, C54A, C54R, C55A, C55R, C56A, C56R,
  C57A, C57R, C60A, C60R, CA2_, CA3_, CA4_, CA5_, CA6_, CAD1, CAD2, CAD3,
  CAD4, CAD5, CAD6, CAG, CBG, CCH05, CCH06, CCH07, CCH10, CCH11, CCH12,
  CCH13, CCH14, CCH33, CCH34, CCH35, CCHG_, CCS0, CCS0_, CDUCLK, CDUSTB_,
  CDUXD, CDUXDM, CDUXDP, CDUYD, CDUYDM, CDUYDP, CDUZD, CDUZDM, CDUZDP,
  CEBG, CFBG, CG11, CG12, CG13, CG14, CG15, CG16, CG21, CG22, CG23, CG24,
  CG26, CGCWAR, CGG, CGMC, CH01, CH02, CH03, CH04, CH05, CH06, CH07, CH0705,
  CH0706, CH0707, CH08, CH09, CH10, CH11, CH1108, CH1109, CH1110, CH1111,
  CH1112, CH1113, CH1114, CH1116, CH12, CH1207, CH1208, CH1209, CH1210,
  CH1211, CH1212, CH1213, CH1214, CH1216, CH13, CH1301, CH1302, CH1303,
  CH1304, CH1305, CH1306, CH1307, CH1308, CH1309, CH1310, CH1311, CH1316,
  CH14, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406, CH1407, CH1408,
  CH1409, CH1410, CH1411, CH1412, CH1413, CH1414, CH1416, CH1501, CH1502,
  CH1503, CH1504, CH1505, CH16, CH1601, CH1602, CH1603, CH1604, CH1605,
  CH1606, CH1607, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207,
  CH3208, CH3209, CH3210, CH3310, CH3311, CH3312, CH3313, CH3314, CH3316,
  CHAT01, CHAT02, CHAT03, CHAT04, CHAT05, CHAT06, CHAT07, CHAT08, CHAT09,
  CHAT10, CHAT11, CHAT12, CHAT13, CHAT14, CHBT01, CHBT02, CHBT03, CHBT04,
  CHBT05, CHBT06, CHBT07, CHBT08, CHBT09, CHBT10, CHBT11, CHBT12, CHBT13,
  CHBT14, CHINC, CHINC_, CHOR01_, CHOR02_, CHOR03_, CHOR04_, CHOR05_, CHOR06_,
  CHOR07_, CHOR08_, CHOR09_, CHOR10_, CHOR11_, CHOR12_, CHOR13_, CHOR14_,
  CHOR16_, CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_,
  CHWL08_, CHWL09_, CHWL10_, CHWL11_, CHWL12_, CHWL13_, CHWL14_, CHWL16_,
  CI, CI01_, CI02_, CI03_, CI04_, CI05_, CI06_, CI07_, CI08_, CI09_, CI10_,
  CI11_, CI12_, CI13_, CI14_, CI15_, CI16_, CIFF, CINORM, CI_, CKTAL_,
  CLEARA, CLEARB, CLEARC, CLEARD, CLG1G, CLG2G, CLK, CLROPE, CLXC, CNTOF9,
  CNTRSB_, CO02, CO04, CO06, CO08, CO10, CO12, CO14, CO16, COARSE, COMACT,
  CON1, CON2, CON3, CQG, CSG, CSQG, CT, CTPLS_, CTROR, CTROR_, CT_, CUG,
  CXB0_, CXB1_, CXB2_, CXB3_, CXB4_, CXB5_, CXB6_, CXB7_, CYL_, CYR_, CZG,
  DAS0, DAS0_, DAS1, DAS1_, DATA_, DBLTST, DCA0, DCS0, DIM0, DIM0_, DINC,
  DINCNC_, DINC_, DISDAC, DIVSTG, DIV_, DKCTR1, DKCTR1_, DKCTR2, DKCTR2_,
  DKCTR3, DKCTR3_, DKCTR4, DKCTR4_, DKCTR5, DKCTR5_, DKDATA, DKDATB, DKDAT_,
  DLKCLR, DLKPLS, DLKRPT, DNRPTA, DOFILT, DOSCAL, DRPRST, DV0, DV0_, DV1,
  DV1376, DV1376_, DV1B1B, DV1_, DV376, DV3764, DV376_, DV4, DV4B1B, DV4_,
  DVST, DVST_, DVXP1, DXCH0, E5, E6, E7_, EAC_, EAD09, EAD09_, EAD10, EAD10_,
  EAD11, EAD11_, EB10, EB10_, EB11, EB11_, EB9, EB9_, EDOP_, EDSET, ELSNCM,
  ELSNCN, EMSD, EMSm, EMSp, END, ENERIM, ENEROP, ERAS, ERAS_, ERRST, EVNSET,
  EVNSET_, EXST0_, EXST1_, EXT, EXTPLS, F01A, F01B, F01C, F01D, F02A, F02B,
  F03A, F03B, F03B_, F04A, F04B, F04B_, F05A, F05A_, F05B, F05B_, F05D,
  F06A, F06B, F06B_, F07A, F07A_, F07B, F07B_, F07C_, F07D_, F08A, F08B,
  F08B_, F09A, F09A_, F09B, F09B_, F09D, F10A, F10AS0, F10A_, F10B, F10B_,
  F11, F11A, F11B, F11_, F12, F12A, F12B, F12B_, F12_, F13, F13A, F13B,
  F13_, F14, F14A, F14B, F14H, F14_, F15, F15A, F15B, F15_, F16, F16A,
  F16B, F16_, F17A, F17A_, F17B, F17B_, F18A, F18AX, F18A_, F18B, F18B_,
  F19A, F19B, F20A, F20B, F21A, F21B, F22A, F22B, F23A, F23B, F24A, F24B,
  F25A, F25B, F26A, F26B, F27A, F27B, F28A, F28B, F29A, F29B, F30A, F30B,
  F31A, F31B, F32A, F32B, F33A, F33B, F5ASB0, F5ASB0_, F5ASB2, F5ASB2_,
  F5BSB2, F5BSB2_, F7CSB1_, FB11, FB11_, FB12, FB12_, FB13, FB13_, FB14,
  FB14_, FB16, FB16_, FETCH0, FETCH0_, FETCH1, FF1109, FF1109_, FF1110,
  FF1110_, FF1111, FF1111_, FF1112, FF1112_, FILTIN, FLASH, FLASH_, FNERAS_,
  FS01, FS01_, FS02, FS02A, FS03, FS03A, FS04, FS04A, FS05, FS05A, FS05_,
  FS06, FS06_, FS07, FS07A, FS07_, FS08, FS08_, FS09, FS09_, FS10, FS11,
  FS12, FS13, FS13_, FS14, FS15, FS16, FS17, FS18, FS19, FS20, FS21, FS22,
  FS23, FS24, FS25, FS26, FS27, FS28, FS29, FS30, FS31, FS32, FS33, FUTEXT,
  G01, G01A, G01A_, G01ED, G01_, G02, G02ED, G02_, G03, G03ED, G03_, G04,
  G04ED, G04_, G05, G05ED, G05_, G06, G06ED, G06_, G07, G07ED, G07_, G08,
  G08_, G09, G09_, G10, G10_, G11, G11_, G12, G12_, G13, G13_, G14, G14_,
  G15, G15_, G16, G16A_, G16SW_, G16_, G2LSG, G2LSG_, GEM01, GEM02, GEM03,
  GEM04, GEM05, GEM06, GEM07, GEM08, GEM09, GEM10, GEM11, GEM12, GEM13,
  GEM14, GEM16, GEMP, GEQZRO_, GINH, GNHNC, GNZRO, GOJ1, GOJ1_, GOJAM,
  GOJAM_, GOSET_, GTONE, GTRST, GTRST_, GTSET, GTSET_, GYENAB, GYROD, GYRRST,
  GYRSET, GYXM, GYXP, GYYM, GYYP, GYZM, GYZP, HERB, HIGH0_, HIGH1_, HIGH2_,
  HIGH3_, HIMOD, HNDRPT, IC1, IC10, IC10_, IC11, IC11_, IC12, IC12_, IC13,
  IC13_, IC14, IC15, IC15_, IC16, IC16_, IC17, IC2, IC2_, IC3, IC3_, IC4,
  IC4_, IC5, IC5_, IC6, IC7, IC8_, IC9, IC9_, IHENV, IIP, IIP_, IL01, IL01_,
  IL02, IL02_, IL03, IL03_, IL04, IL04_, IL05, IL05_, IL06, IL06_, IL07,
  IL07_, ILP, ILP_, INCR0, INCSET_, INHINT, INHPLS, INKBT1, INKL, INKL_,
  INLNKM, INLNKP, INOTLD, INOTRD, INOUT, INOUT_, ISSTDC, ISSWAR, KRPT,
  KRPTA_, KY1RST, KY2RST, KYRLS, KYRPT1, KYRPT2, L01_, L02A_, L02_, L03_,
  L04_, L05_, L06_, L07_, L08_, L09_, L10_, L11_, L12_, L13_, L14_, L15A_,
  L15_, L16_, L2GDG_, L2GD_, LOMOD, LOW0_, LOW1_, LOW2_, LOW3_, LOW4_,
  LOW5_, LOW6_, LOW7_, LRRANG, LRRST, LRSYNC, LRXVEL, LRYVEL, LRZVEL, LXCH0,
  MAMU, MASK0, MASK0_, MBR1, MBR2, MCDU, MCDU_, MCRO_, MCTRAL_, MDT01,
  MDT02, MDT03, MDT04, MDT05, MDT06, MDT07, MDT08, MDT09, MDT10, MDT11,
  MDT12, MDT13, MDT14, MDT15, MDT16, MGOJAM, MGP_, MIIP, MINC, MINC_, MINHL,
  MINKL, MISSX, MISSY, MISSZ, MKRPT, MLDCH, MLOAD, MNHNC, MNHRPT, MNHSBF,
  MNISQ, MON800, MONEX, MONEX_, MONPAR, MONWBK, MONWT, MON_, MONpCH, MOSCAL_,
  MOUT, MOUT_, MP0, MP0T10, MP0_, MP1, MP1_, MP3, MP3A, MP3_, MPAL_, MPIPAL_,
  MRAG, MRCH, MRDCH, MREAD, MREQIN, MRGG, MRLG, MROLGT, MRPTAL_, MRSC,
  MRULOG, MSBSTP, MSCAFL_, MSCDBL_, MSP, MSQ10, MSQ11, MSQ12, MSQ13, MSQ14,
  MSQ16, MSQEXT, MST1, MST2, MST3, MSTP, MSTPIT_, MSTRT, MSTRTP, MSU0,
  MSU0_, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11,
  MT12, MTCAL_, MTCSAI, MTCSA_, MVFAIL_, MWAG, MWARNF_, MWATCH_, MWBBEG,
  MWBG, MWCH, MWEBG, MWFBG, MWG, MWL01, MWL02, MWL03, MWL04, MWL05, MWL06,
  MWL07, MWL08, MWL09, MWL10, MWL11, MWL12, MWL13, MWL14, MWL15, MWL16,
  MWLG, MWQG, MWSG, MWYG, MWZG, NDR100_, NDX0, NDX0_, NDXX1, NDXX1_, NEAC,
  NEXST0, NEXST0_, NHALGA, NISQ, NISQL_, NISQ_, NOTEST, NOTEST_, NOXM,
  NOXP, NOYM, NOYP, NOZM, NOZP, OCTAD2, OCTAD3, OCTAD4, OCTAD5, OCTAD6,
  ODDSET_, ONE, OPEROR, ORDRBT, OSCALM, OT1108, OT1110, OT1111, OT1112,
  OT1113, OT1114, OT1116, OT1207, OT1207_, OTLNK0, OTLNK1, OTLNKM, OUTCOM,
  OVF, OVFSTB_, OVF_, OVNHRP, P01, P01_, P02, P02_, P03, P03_, P04, P04A,
  P04_, P05, P05_, PA03, PA03_, PA06, PA06_, PA09, PA09_, PA12, PA12_,
  PA15, PA15_, PALE, PARTC, PB09, PB09_, PB15, PB15_, PC15, PC15_, PCDU,
  PCDU_, PHS2, PHS2_, PHS3_, PHS4, PHS4_, PIFL_, PINC, PINC_, PIPAFL, PIPASW,
  PIPAXm_, PIPAXp_, PIPAYm_, PIPAYp_, PIPAZm_, PIPAZp_, PIPDAT, PIPGXm,
  PIPGXp, PIPGYm, PIPGYp, PIPGZm, PIPGZp, PIPINT, PIPPLS_, PIPSAM, PIPSAM_,
  PIPXM, PIPXP, PIPYM, PIPYP, PIPZM, PIPZP, PONEX, POUT, POUT_, PRINC,
  PRPOR1, PRPOR2, PRPOR3, PRPOR4, PSEUDO, PTWOX, Q2A, QC0, QC0_, QC1_,
  QC2_, QC3_, QXCH0, QXCH0_, R15, R1C, R1C_, R6, RAD, RADRG, RADRPT, RADRZ,
  RAG_, RAND0, RA_, RB1, RB1F, RB1_, RB2, RBBEG_, RBBK, RBHG_, RBLG_, RBSQ,
  RB_, RCG_, RCH05_, RCH06_, RCH07_, RCH10_, RCH11_, RCH12_, RCH13_, RCH14_,
  RCH15_, RCH16_, RCH30_, RCH31_, RCH32_, RCH33_, RCHAT_, RCHBT_, RCHG_,
  RCH_, RC_, RCmXmP, RCmXmY, RCmXpP, RCmXpY, RCmYmR, RCmYpR, RCmZmR, RCmZpR,
  RCpXmP, RCpXmY, RCpXpP, RCpXpY, RCpYmR, RCpYpR, RCpZmR, RCpZpR, RDBANK,
  RDOUT_, READ0, READ0_, REBG_, REDRST, RELPLS, RESETA, RESETB, RESETC,
  RESETD, RESTRT, REX, REY, RFBG_, RGG1, RGG_, RG_, RHCGO, RILP1, RILP1_,
  RINGA_, RINGB_, RL01_, RL02_, RL03_, RL04_, RL05_, RL06_, RL07_, RL08_,
  RL09_, RL10BB, RL10_, RL11_, RL12_, RL13_, RL14_, RL15_, RL16, RL16_,
  RLG1, RLG2, RLG3, RLG_, RLYB01, RLYB02, RLYB03, RLYB04, RLYB05, RLYB06,
  RLYB07, RLYB08, RLYB09, RLYB10, RLYB11, RL_, RNRADM, RNRADP, ROPER, ROPES,
  ROPET, ROP_, ROR0, RPTA12, RPTAD3, RPTAD4, RPTAD5, RPTAD6, RPTFRC, RPTSET,
  RQ, RQG_, RQ_, RRPA, RRPA1_, RRRANG, RRRARA, RRRST, RRSYNC, RSCG_, RSCT,
  RSCT_, RSC_, RSM3, RSM3_, RSSB, RSTKX_, RSTKY_, RSTK_, RSTRT, RSTSTG,
  RT, RT_, RUG_, RULOG_, RUPT0, RUPT0_, RUPT1, RUPT1_, RUPTOR_, RUSG_,
  RUS_, RU_, RXOR0, RXOR0_, RYWD12, RYWD13, RYWD14, RYWD16, RZG_, RZ_,
  S01, S01_, S02, S02_, S03, S03_, S04, S04_, S05, S05_, S06, S06_, S07,
  S07_, S08, S08A, S08A_, S08_, S09, S09_, S10, S10_, S11, S11_, S12, S12_,
  S4BOFF, S4BSEQ, S4BTAK, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08,
  SA09, SA10, SA11, SA12, SA13, SA14, SA16, SAP, SB0, SB0_, SB1, SB1_,
  SB2, SB2_, SB4, SBE, SBESET, SBF, SBFSET, SBY, SBYEXT, SBYLIT, SBYREL_,
  SCAD, SCADBL, SCAD_, SCAS10, SCAS17, SETAB, SETAB_, SETCD, SETCD_, SETEK,
  SGUM, SH3MS_, SHAFTD, SHANC, SHANC_, SHFTDM, SHFTDP, SHIFT, SHIFT_, SHINC,
  SHINC_, SQ0_, SQ1_, SQ2_, SQ3_, SQ4_, SQ5, SQ5QC0_, SQ5_, SQ6_, SQ7_,
  SQEXT, SQEXT_, SQR10, SQR10_, SQR11, SQR12, SQR12_, SQR13, SQR14, SQR16,
  SR_, ST0_, ST1, ST1376_, ST1D, ST1_, ST2, ST2_, ST376, ST376_, ST3_,
  ST4_, STARON, STBE, STBF, STD2, STFET1_, STG1, STG2, STG3, STNDBY, STNDBY_,
  STOP, STOPA, STOP_, STORE1, STORE1_, STR14, STR19, STR210, STR311, STR412,
  STR58, STR912, STRGAT, STRT1, STRTFC, SU0, SUMA01_, SUMA02_, SUMA03_,
  SUMA04_, SUMA05_, SUMA06_, SUMA07_, SUMA08_, SUMA09_, SUMA10_, SUMA11_,
  SUMA12_, SUMA13_, SUMA14_, SUMA15_, SUMA16_, SUMB01_, SUMB02_, SUMB03_,
  SUMB04_, SUMB05_, SUMB06_, SUMB07_, SUMB08_, SUMB09_, SUMB10_, SUMB11_,
  SUMB12_, SUMB13_, SUMB14_, SUMB15_, SUMB16_, SYNC14_, SYNC4_, T01, T01DC_,
  T01_, T02, T02DC_, T02_, T03, T03DC_, T03_, T04, T04_, T05, T05_, T06,
  T06DC_, T06_, T07, T07DC_, T07_, T08, T08DC_, T08_, T09, T09DC_, T09_,
  T10, T10DC_, T10_, T11, T11_, T12, T12A, T12DC_, T12SET, T12USE_, T12_,
  T1P, T2P, T3P, T4P, T5P, T6ON_, T6P, T6RPT, T7PHS4, T7PHS4_, TC0, TC0_,
  TCF0, TCSAJ3, TCSAJ3_, TEMPIN_, THRSTD, THRSTm, THRSTp, TIMR, TL15, TMPCAU,
  TMPOUT, TMZ_, TOV_, TPARG_, TPGE, TPGF, TPORA_, TPOR_, TPZG_, TRNDM,
  TRNDP, TRP31A, TRP31B, TRP32, TRSM, TRSM_, TRUND, TS0, TS0_, TSGN2, TSGN_,
  TSGU_, TSUDO_, TT_, TVCNAB, TWOX, U2BBK, U2BBKG_, UNF, UNF_, UPL0_, UPL1_,
  UPLACT, UPRUPT, US2SG, VNFLSH, W1110, WAG_, WALSG, WALSG_, WAND0, WARN,
  WATCH, WATCHP, WATCH_, WA_, WBBEG_, WBG_, WB_, WCH05_, WCH06_, WCH07_,
  WCH10_, WCH11_, WCH12_, WCH13_, WCH14_, WCH34_, WCH35_, WCHG_, WCH_,
  WDORDR, WEBG_, WEDOPG_, WEX, WEY, WFBG_, WG1G_, WG2G_, WG3G_, WG4G_,
  WG5G_, WGA_, WGNORM, WG_, WHOMP, WHOMPA, WHOMP_, WL01, WL01_, WL02, WL02_,
  WL03, WL03_, WL04, WL04_, WL05, WL05_, WL06, WL06_, WL07, WL07_, WL08,
  WL08_, WL09, WL09_, WL10, WL10_, WL11, WL11_, WL12, WL12_, WL13, WL13_,
  WL14, WL14_, WL15, WL15_, WL16, WL16_, WLG_, WL_, WOR0, WOR0_, WOVR,
  WOVR_, WQG_, WQ_, WRD1B1, WRD1BP, WRD2B2, WRD2B3, WRITE0, WRITE0_, WSCG_,
  WSC_, WSG_, WSQG_, WS_, WT, WT_, WY12_, WYDG_, WYDLOG_, WYD_, WYHIG_,
  WYLOG_, WY_, WZG_, WZ_, XB0, XB0E, XB0_, XB1, XB1E, XB1_, XB2, XB2E,
  XB2_, XB3, XB3E, XB3_, XB4, XB4E, XB4_, XB5, XB5E, XB5_, XB6, XB6E, XB6_,
  XB7, XB7E, XB7_, XLNK0_, XLNK1_, XT0, XT0E, XT0_, XT1, XT1E, XT1_, XT2,
  XT2E, XT2_, XT3, XT3E, XT3_, XT4, XT4E, XT4_, XT5, XT5E, XT5_, XT6, XT6E,
  XT6_, XT7, XT7E, XT7_, XUY01_, XUY02_, XUY03_, XUY04_, XUY05_, XUY06_,
  XUY07_, XUY08_, XUY09_, XUY10_, XUY11_, XUY12_, XUY13_, XUY14_, XUY15_,
  XUY16_, YB0, YB0E, YB0_, YB1, YB1E, YB1_, YB2, YB2E, YB2_, YB3, YB3E,
  YB3_, YT0, YT0E, YT0_, YT1, YT1E, YT1_, YT2, YT2E, YT2_, YT3, YT3E, YT3_,
  YT4, YT4E, YT4_, YT5, YT5E, YT5_, YT6, YT6E, YT6_, YT7, YT7E, YT7_, Z01_,
  Z02_, Z03_, Z04_, Z05_, Z06_, Z07_, Z08_, Z09_, Z10_, Z11_, Z12_, Z13_,
  Z14_, Z15_, Z16_, ZAP, ZAP_, ZEROPT, ZID, ZIMCDU, ZIP, ZIPCI, ZOPCDU,
  ZOUT, ZOUT_, d10XP1, d10XP6, d10XP8, d11XP2, d12KPPS, d16CNT, d1CNT,
  d1XP10, d25KPPS, d2PP1, d2XP3, d2XP5, d2XP7, d2XP8, d30SUM, d32004K,
  d3200A, d3200B, d3200C, d3200D, d32CNT, d3XP2, d3XP6, d3XP7, d4XP11,
  d4XP5, d50SUM, d5XP11, d5XP12, d5XP15, d5XP21, d5XP28, d5XP4, d6XP5,
  d6XP8, d7XP14, d7XP19, d7XP4, d7XP9, d800RST, d800SET, d8PP4, d8XP5,
  d8XP6, d9XP1, d9XP5;

A1 iA1 (
  rst, CGA1, FS01_, RCHAT_, RCHBT_, F03B, F07A, F09A, F17A, F18A, F18A_,
  F25A, FS06, FS07, FS07_, FS08, CHAT01, CHAT02, CHAT03, CHAT04, CHAT05,
  CHAT06, CHAT07, CHAT08, CHAT09, CHAT10, CHAT11, CHAT12, CHAT13, CHAT14,
  CHBT01, CHBT02, CHBT03, CHBT04, CHBT05, CHBT06, CHBT07, CHBT08, CHBT09,
  CHBT10, CHBT11, CHBT12, CHBT13, CHBT14, F02A, F02B, F03A, F03B_, F04A,
  F04B, F05A, F05B, F06A, F06B, F07A_, F07B, F08A, F08B, F09B, F10A, F10B,
  F11A, F11B, F12A, F12B, F13A, F13B, F14A, F14B, F15A, F15B, F16A, F16B,
  F17B, F18AX, F18B, F19A, F19B, F20A, F20B, F21A, F21B, F22A, F22B, F23A,
  F23B, F24A, F24B, F25B, F26A, F26B, F27A, F27B, F28A, F28B, F29A, F29B,
  F30A, F30B, F31A, F31B, F32A, F32B, F33A, F33B, FS02, FS02A, FS03, FS03A,
  FS04, FS04A, FS05, FS05A, FS06_, FS07A, FS08_, FS09, FS10, FS11, FS12,
  FS13, FS14, FS15, FS16, FS17, FS18, FS19, FS20, FS21, FS22, FS23, FS24,
  FS25, FS26, FS27, FS28, FS29, FS30, FS31, FS32, FS33
);
defparam iA1.GATE_DELAY = GATE_DELAY;

A2 iA2 (
  rst, ALGA, CGA2, CLOCK, GOJ1, MP3A, MSTP, MSTRTP, SBY, STRT1, STRT2, WL15,
  WL15_, WL16, WL16_, CINORM, EVNSET, EVNSET_, GOJAM, GOJAM_, MGOJAM, MONWT,
  MSTPIT_, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11,
  MT12, ODDSET_, OVFSTB_, P01_, P02, P02_, P03, P03_, P04, P05, P05_, PHS4,
  PHS4_, Q2A, RINGA_, RINGB_, RT, STOP, STOPA, T02, T02DC_, T03, T03DC_,
  T06, T06DC_, T08, T08DC_, T10, T10DC_, T12DC_, WT, WT_, CLK, CT, CT_, EDSET,
  F01A, F01B, F01C, F01D, FS01, FS01_, GOSET_, OVF, OVF_, P01, P04_, PHS2,
  PHS2_, RT_, SB0, SB1, SB2, SB4, STOP_, T01, T01DC_, T01_, T02_, T03_, T04,
  T04_, T05, T05_, T06_, T07, T07DC_, T07_, T08_, T09, T09DC_, T09_, T10_,
  T11, T11_, T12, T12SET, T12_, TT_, UNF, UNF_
);
defparam iA2.GATE_DELAY = GATE_DELAY;

A3 iA3 (
  rst, BR1B2B, BR2_, CGA3, CT_, DBLTST, EXT, EXTPLS, FS09, FS10, GOJAM, INHPLS,
  INKL, KRPT, MNHRPT, MTCSAI, NISQ, ODDSET_, OVNHRP, PHS2_, RELPLS, RT_,
  RUPTOR_, RXOR0, ST0_, ST1_, ST3_, STD2, T01_, T02, T07DC_, T12_, WL10_,
  WL11_, WL12_, WL13_, WL14_, WL16_, WT_, d5XP4, CON1, CON2, EXST0_, INKBT1,
  MIIP, MINHL, MSQ10, MSQ11, MSQ12, MSQ13, MSQ14, MSQ16, MSQEXT, MTCSA_,
  NEXST0, QC0, QC0_, QC1_, QC2_, QC3_, RPTSET, SCAS10, SQ0_, SQ1_, SQ2_,
  SQ3_, SQ4_, SQ5, SQ6_, SQ7_, SQEXT, SQEXT_, T07, TCSAJ3, TS0, AD0, ADS0,
  AUG0, AUG0_, BMF0, BMF0_, BZF0, BZF0_, CCS0, CCS0_, CSQG, DAS0, DAS0_,
  DAS1, DAS1_, DCA0, DCS0, DIM0, DIM0_, DXCH0, EXST1_, FUTEXT, GOJ1, GOJ1_,
  IC1, IC10, IC10_, IC11, IC12, IC12_, IC13, IC13_, IC14, IC15, IC15_, IC16,
  IC16_, IC17, IC2, IC2_, IC3, IC3_, IC4, IC4_, IC5, IC5_, IC6, IC7, IC8_,
  IC9, IC9_, IIP, IIP_, INCR0, INHINT, LXCH0, MASK0, MASK0_, MP0, MP0_, MP1,
  MP1_, MP3, MP3_, MSU0, MSU0_, NDX0, NDX0_, NDXX1, NDXX1_, NEXST0_, NISQL_,
  QXCH0, QXCH0_, RBSQ, RPTFRC, RSM3, RSM3_, SQ5QC0_, SQ5_, SQR10, SQR10_,
  SQR11, SQR12, SQR12_, SQR13, SQR14, SQR16, STRTFC, SU0, TC0, TC0_, TCF0,
  TCSAJ3_, TS0_, WSQG_
);
defparam iA3.GATE_DELAY = GATE_DELAY;

A4 iA4 (
  rst, CGA4, DVST, EXST0_, EXST1_, GEQZRO_, GOJAM, IC12, IC13, INKL, L15_,
  MP0_, MP1, MP3_, MTCSAI, NDR100_, OVF_, PHS2_, PHS3_, PHS4, PHS4_, QC0_,
  QC1_, QC2_, QC3_, RSM3, RSM3_, RSTSTG, SQ0_, SQ1_, SQ2_, SQEXT, SQEXT_,
  SQR10, SQR10_, SQR12_, ST1, ST2, STORE1_, STRTFC, SUMA16_, SUMB16_, T01,
  T01_, T02_, T03_, T04_, T05_, T06_, T07_, T08_, T09_, T10_, T11_, T12_,
  TOV_, TPZG_, TRSM, TS0_, TSGU_, UNF_, WL01_, WL02_, WL03_, WL04_, WL05_,
  WL06_, WL07_, WL08_, WL09_, WL10_, WL11_, WL12_, WL13_, WL14_, WL15_, WL16_,
  XB7_, XT1_, d7XP14, BR1, BR1_, BR2, BR2_, CI_, DV0_, DV1_, DV4, DVST_,
  L16_, MBR1, MBR2, MP3A, MRSC, MST1, MST2, MST3, R1C_, RA_, RB1_, RB_, RC_,
  ST0_, TL15, TMZ_, TRSM_, TSGN2, TSGN_, WG_, WL_, WY_, d2PP1, B15X, BR12B,
  BR12B_, BR1B2, BR1B2B, BR1B2B_, BR1B2_, BRDIF_, DIVSTG, DIV_, DV0, DV1,
  DV1376, DV1376_, DV376, DV3764, DV376_, DV4_, INOUT, INOUT_, KRPT, MP0T10,
  PRINC, R15, RAND0, RB2, READ0, READ0_, ROR0, RRPA, RSC_, RUPT0, RUPT0_,
  RUPT1, RUPT1_, RXOR0, RXOR0_, SGUM, ST1376_, ST1D, ST1_, ST376, ST376_,
  ST3_, ST4_, STD2, STG1, STG2, STG3, T12USE_, WAND0, WCH_, WOR0, WOR0_,
  WRITE0, WRITE0_, d1XP10, d2XP3, d2XP5, d3XP2, d3XP7, d4XP11, d4XP5, d5XP11,
  d5XP28, d5XP4, d6XP5, d7XP19, d8PP4, d8XP5, d8XP6, d9XP1
);
defparam iA4.GATE_DELAY = GATE_DELAY;

A5 iA5 (
  rst, ADS0, BR1, BR12B_, BR1B2_, BR1_, BR2, BR2_, BRDIF_, C24A, C25A, C26A,
  C27A, C30A, C37P, C40P, C41P, C42P, C43P, C44P, CCS0, CCS0_, CGA5, CHINC_,
  DAS0, DAS0_, DAS1, DAS1_, DIV_, DV1, DV1_, DV4, DV4_, DXCH0, EDSET, FETCH0,
  FETCH0_, GOJ1, GOJ1_, GOJAM, IC1, IC10, IC10_, IC11_, IC12, IC12_, IC13,
  IC14, IC15_, IC16, IC16_, IC2, IC2_, IC3, IC4, IC5, IC5_, IC8_, IC9, INCSET_,
  INKL_, INOUT, INOUT_, MASK0, MASK0_, MONWBK, MONpCH, MP0, MP3, MP3_, MSU0,
  MSU0_, NDX0_, PRINC, QXCH0_, RAND0, READ0, ROR0, RSM3, RSM3_, RUPT0, RXOR0,
  RXOR0_, S11, S12, SHANC_, SHIFT, SHIFT_, STD2, STFET1_, T01, T01_, T02_,
  T03_, T04_, T05_, T06_, T07_, T08_, T09_, T10_, T11_, T12, T12USE_, T12_,
  TC0, TC0_, TCF0, TCSAJ3_, TS0, TS0_, WAND0, WOR0, XT0_, XT2_, XT3_, XT4_,
  XT5_, XT6_, YB0_, YT0_, d4XP5, d5XP11, A2X_, CI_, DV1B1B, MONEX_, P03,
  PARTC, RA_, RB_, RC_, RG_, RL_, RU_, RZ_, ST2_, TMZ_, TOV_, TSGN_, WA_,
  WB_, WG_, WL_, WS_, WY12_, WYD_, WY_, WZ_, Z15_, Z16_, d10XP6, DV4B1B,
  DVST, GNHNC, NDR100_, NISQ_, OCTAD2, OCTAD3, OCTAD4, OCTAD5, OCTAD6, PINC,
  PINC_, PTWOX, R6, RAD, RL10BB, RQ, RSCT, RSTRT, RSTSTG, SCAD, SCAD_, TPZG_,
  TRSM, TSUDO_, U2BBK, d10XP1, d10XP8, d11XP2, d2XP7, d2XP8, d3XP6, d5XP12,
  d5XP15, d5XP21, d6XP8, d7XP4, d7XP9, d9XP5
);
defparam iA5.GATE_DELAY = GATE_DELAY;

A6 iA6 (
  rst, AD0, ADS0, AUG0_, B15X, BR1, BR12B_, BR1B2B, BR1B2B_, BR1B2_, BR1_,
  BR2_, CCS0, CCS0_, CDUSTB_, CGA6, DAS0, DAS1, DAS1_, DCA0, DCS0, DIM0_,
  DINC, DINC_, DIVSTG, DV0, DV1376, DV1376_, DV376_, DV4B1B, DV4_, DXCH0,
  FETCH1, GOJAM, IC11, IC15, IC17, IC6, IC7, IC9, INCR0, INKL, INOTLD, L01_,
  L02A_, L15A_, MASK0, MCDU, MINC, MON_, MONpCH, MP0T10, MP1, MP1_, MP3_,
  MSU0, NDXX1_, P01, P04, P05_, PCDU, PHS4_, PINC, PRINC, PTWOX, R15, R6,
  RADRG, RADRZ, RAND0, RBSQ, RRPA, RSTK_, RUPT0, RUPT1, S01, S01_, S02, S02_,
  S03, S03_, S04, S04_, S05, S05_, S06, S06_, S07, S07_, SHIFT, STBE, STBF,
  STFET1_, STOP_, STRT2, SU0, T01, T01_, T02, T02_, T03, T03_, T04, T04_,
  T05, T06, T06_, T07, T07_, T08, T08_, T09, T10, T10_, T11, T11_, T12, T12USE_,
  TL15, WAND0, d10XP1, d10XP8, d11XP2, d1XP10, d2XP3, d2XP5, d2XP7, d2XP8,
  d3XP2, d3XP6, d3XP7, d4XP11, d5XP12, d5XP15, d5XP21, d5XP28, d5XP4, d6XP5,
  d6XP8, d7XP19, d7XP4, d7XP9, d8PP4, d8XP6, d9XP1, d9XP5, IL01, IL01_, IL02,
  IL02_, IL03, IL03_, IL04, IL04_, IL05, IL05_, IL06, IL06_, IL07, IL07_,
  MONEX_, RB_, RC_, RDBANK, RPTSET, RSTKX_, RSTKY_, RU_, ST2_, WG_, WSC_,
  WY_, ZIPCI, d2PP1, A2X_, BXVX, CGMC, CI_, CLXC, DVXP1, EXT, L2GD_, MCRO_,
  MONEX, MOUT, NEAC, PIFL_, PONEX, POUT, PSEUDO, R1C_, RB1F, RB1_, RCH_,
  RG_, RUS_, RZ_, ST1, ST2, TIMR, TOV_, TSGU_, TWOX, WA_, WB_, WL_, WOVR,
  WQ_, WS_, WYD_, WZ_, ZAP, ZAP_, ZIP, ZOUT, d7XP14
);
defparam iA6.GATE_DELAY = GATE_DELAY;

A7 iA7 (
  rst, A2X_, CGA7, CGMC, CI, CT_, CYL_, CYR_, EAC_, EAD09, EAD09_, EAD10,
  EAD10_, EAD11, EAD11_, EDOP_, GINH, L15_, L2GD_, NEAC, P04_, PIFL_, PIPPLS_,
  RA_, RB_, RCHG_, RC_, RG_, RL10BB, RL_, RQ_, RSCG_, RT_, RUS_, RU_, RZ_,
  SB2_, SHIFT, SR_, STFET1_, T10_, TT_, U2BBK, WA_, WB_, WCHG_, WGA_, WG_,
  WL_, WQ_, WSCG_, WS_, WT_, WY12_, WYD_, WY_, WZ_, XB0_, XB1_, XB2_, XB3_,
  XB4_, XB5_, XB6_, XT0_, ZAP_, CIFF, CINORM, CSG, CUG, G2LSG, MRAG, MRGG,
  MRLG, MRULOG, MWAG, MWBBEG, MWBG, MWEBG, MWFBG, MWG, MWLG, MWQG, MWSG,
  MWYG, MWZG, P04A, RBBK, RGG1, RGG_, RLG1, RLG2, RLG3, RLG_, WALSG, WSG_,
  YT0E, YT1E, YT2E, YT3E, YT4E, YT5E, YT6E, YT7E, A2XG_, CAG, CBG, CEBG,
  CFBG, CGG, CI01_, CLG1G, CLG2G, CQG, CZG, G2LSG_, L2GDG_, PIPSAM, RAG_,
  RBBEG_, RBHG_, RBLG_, RCG_, REBG_, RFBG_, RQG_, RUG_, RULOG_, RUSG_, RZG_,
  WAG_, WALSG_, WBBEG_, WBG_, WEBG_, WEDOPG_, WFBG_, WG1G_, WG2G_, WG3G_,
  WG4G_, WG5G_, WGNORM, WLG_, WQG_, WYDG_, WYDLOG_, WYHIG_, WYLOG_, WZG_,
  YT0, YT0_, YT1, YT1_, YT2, YT2_, YT3, YT3_, YT4, YT4_, YT5, YT5_, YT6,
  YT6_, YT7, YT7_
);
defparam iA7.GATE_DELAY = GATE_DELAY;

A8 iA8 (
  rst, A2XG_, CAG, CBG, CGA8, CGG, CH01, CH02, CH03, CH04, CI01_, CLG1G,
  CLXC, CQG, CUG, CZG, G01ED, G02ED, G03ED, G04ED, G05ED, G06ED, G07_, G2LSG_,
  L2GDG_, MCRO_, MDT01, MDT02, MDT03, MDT04, MONEX, PONEX, R15, R1C, RAG_,
  RB1, RB2, RBLG_, RCG_, RGG_, RLG_, RQG_, RULOG_, RZG_, S08, S08_, SA01,
  SA02, SA03, SA04, SETAB_, SETCD_, TWOX, WAG_, WALSG_, WBG_, WG1G_, WG3G_,
  WG4G_, WL05_, WL06_, WL16_, WLG_, WQG_, WYDG_, WYDLOG_, WYLOG_, WZG_, XUY05_,
  XUY06_, CI02_, CI03_, CI04_, CO04, CO06, G01_, G02_, G03_, G04_, G05_,
  G06_, GEM01, GEM02, GEM03, GEM04, L01_, L02_, L03_, MWL01, MWL02, MWL03,
  MWL04, RL01_, RL02_, RL03_, RL04_, S08A, S08A_, SUMA04_, WL01_, WL02_,
  WL03_, WL04_, XUY03_, XUY04_, A01_, A02_, A03_, A04_, CI05_, CLEARA, CLEARB,
  CLEARC, CLEARD, G01, G02, G03, G04, L04_, SUMA01_, SUMA02_, SUMA03_, SUMB01_,
  SUMB02_, SUMB03_, SUMB04_, WL01, WL02, WL03, WL04, XUY01_, XUY02_, Z01_,
  Z02_, Z03_, Z04_
);
defparam iA8.GATE_DELAY = GATE_DELAY;

A9 iA9 (
  rst, A2XG_, CAG, CBG, CGA9, CGG, CH05, CH06, CH07, CH08, CI05_, CLG1G,
  CLXC, CO06, CQG, CUG, CZG, G07ED, G09_, G10_, G11_, G2LSG_, L04_, L2GDG_,
  MDT05, MDT06, MDT07, MDT08, MONEX, PIPAXm_, PIPAXp_, PIPAYp_, PIPSAM, R1C,
  RAG_, RBLG_, RCG_, RGG_, RL16_, RLG_, RQG_, RULOG_, RZG_, SA05, SA06, SA07,
  SA08, STRT2, WAG_, WALSG_, WBG_, WG1G_, WG3G_, WG4G_, WL04_, WL09_, WL10_,
  WLG_, WQG_, WYDG_, WYLOG_, WZG_, XUY09_, XUY10_, p4SW, CI06_, CI07_, CI08_,
  CLROPE, CO08, CO10, G05_, G06_, G07_, G08_, GEM05, GEM06, GEM07, GEM08,
  L05_, L06_, L07_, MWL05, MWL06, MWL07, MWL08, PIPSAM_, RL05_, RL06_, ROPER,
  ROPES, ROPET, SUMA07_, WL05_, WL06_, WL07_, WL08_, WL16, XUY07_, XUY08_,
  A05_, A06_, A07_, A08_, CI09_, G05, G06, G07, G08, L08_, PIPGXm, PIPGXp,
  PIPGYp, RL07_, RL08_, SUMA05_, SUMA06_, SUMA08_, SUMB05_, SUMB06_, SUMB07_,
  SUMB08_, WL05, WL06, WL07, WL08, XUY05_, XUY06_, Z05_, Z06_, Z07_, Z08_
);
defparam iA9.GATE_DELAY = GATE_DELAY;

A10 iA10 (
  rst, A2XG_, BK16, CAG, CBG, CGA10, CGG, CH09, CH10, CH11, CH12, CI09_,
  CLG1G, CLXC, CO10, CQG, CUG, CZG, G13_, G14_, G15_, G2LSG_, L08_, L2GDG_,
  MDT09, MDT10, MDT11, MDT12, MONEX, PIPAXm, PIPAXp, PIPAYm_, PIPAYp, PIPAZm_,
  PIPAZp_, PIPSAM_, R1C, RAG_, RBHG_, RBLG_, RCG_, RGG_, RLG_, RQG_, RULOG_,
  RZG_, SA09, SA10, SA11, SA12, WAG_, WALSG_, WBG_, WG1G_, WG3G_, WG4G_,
  WHOMPA, WL08_, WL13_, WL14_, WLG_, WQG_, WYDG_, WYLOG_, WZG_, XUY13_, XUY14_,
  CI10_, CI11_, CI12_, CO04, CO12, CO14, G12_, GEM09, GEM10, GEM11, GEM12,
  L09_, L10_, L11_, MWL09, MWL10, MWL11, MWL12, RL09_, RL10_, RL11_, RL12_,
  RL15_, WL09_, WL10_, WL11_, WL12_, XUY11_, XUY12_, A09_, A10_, A11_, A12_,
  CI13_, G09, G09_, G10, G10_, G11, G11_, G12, L12_, PIPAXm_, PIPAXp_, PIPAYp_,
  PIPGYm, PIPGZm, PIPGZp, SUMA09_, SUMA10_, SUMA11_, SUMA12_, SUMB09_, SUMB10_,
  SUMB11_, SUMB12_, WL09, WL10, WL11, WL12, XUY09_, XUY10_, Z09_, Z10_, Z11_,
  Z12_
);
defparam iA10.GATE_DELAY = GATE_DELAY;

A11 iA11 (
  rst, A2XG_, BXVX, CAG, CBG, CGA11, CGG, CH13, CH14, CH16, CI13_, CLG1G,
  CLG2G, CLXC, CO14, CQG, CUG, CZG, DVXP1, G01_, G16SW_, G2LSG_, GOJAM, GTRST,
  L12_, L2GDG_, MDT13, MDT14, MDT15, MDT16, MONEX, NISQ, ONE, PIPAYm, PIPAZm,
  PIPAZp, R1C, RAG_, RBHG_, RCG_, RGG_, RLG_, RQG_, RUG_, RULOG_, RZG_, SA13,
  SA14, SA16, US2SG, WAG_, WALSG_, WBG_, WG1G_, WG2G_, WG3G_, WG4G_, WG5G_,
  WHOMPA, WL01_, WL02_, WL12_, WLG_, WQG_, WYDG_, WYHIG_, WZG_, XUY01_, XUY02_,
  CI14_, CI15_, CI16_, CO02, CO16, G16_, GEM13, GEM14, GEM16, L13_, L14_,
  L16_, MWL13, MWL14, MWL15, MWL16, RL13_, RL14_, RL15_, RL16, RL16_, SUMA02_,
  SUMA04_, SUMA07_, SUMA12_, SUMA16_, WHOMP, WHOMP_, WL13_, WL14_, WL15_,
  WL16_, XUY15_, XUY16_, Z15_, Z16_, A13_, A14_, A15_, A16_, EAC_, G13, G13_,
  G14, G14_, G15, G15_, G16, GTRST_, L15_, PIPAYm_, PIPAZm_, PIPAZp_, SUMA13_,
  SUMA14_, SUMA15_, SUMB13_, SUMB14_, SUMB15_, SUMB16_, WL13, WL14, WL15,
  WL16, XUY13_, XUY14_, Z13_, Z14_
);
defparam iA11.GATE_DELAY = GATE_DELAY;

A12 iA12 (
  rst, CAD4, CAD5, CAD6, CGA12, CGG, CSG, EB10, EB11_, EB9, G01, G02, G03,
  G04, G05, G06, G07, G08, G09, G10, G11, G12, G13, G14, G15, G16, GOJAM,
  IC15_, L02_, L15_, MONPAR, OCTAD2, R6, RAD, RPTAD4, RPTAD5, RPTAD6, SAP,
  SCAD, SCADBL, SHANC, SHINC, T02_, T03, T04, T05, T07, T10, T12_, T7PHS4_,
  TPARG_, TSUDO_, WEDOPG_, WL01_, WL02_, WL03_, WL04_, WL05_, WL06_, WL07_,
  WL08_, WL09_, WL10_, WL11_, WL12_, WL13_, WL14_, WSG_, XB0_, XB1_, XB2_,
  XB3_, d8XP5, BRXP3, G01A_, GEMP, GNZRO, MGP_, MPAL_, MSCDBL_, MSP, PA03,
  PA03_, PA06, PA06_, PA09, PA09_, PA12, PA12_, PA15, PA15_, RL03_, RL04_,
  RL05_, RL06_, RSC_, S09_, S10_, T03_, T04_, T05_, T07_, T10_, T12A, WG_,
  CYL_, CYR_, EAD09, EAD09_, EAD10, EAD10_, EAD11, EAD11_, EDOP_, EXTPLS,
  G01A, G01ED, G02ED, G03ED, G04ED, G05ED, G06ED, G07ED, G16A_, GEQZRO_,
  GINH, INHPLS, L02A_, L15A_, PALE, PB09, PB09_, PB15, PB15_, PC15, PC15_,
  RADRG, RADRZ, RELPLS, S01, S01_, S02, S02_, S03, S03_, S04, S04_, S05,
  S05_, S06, S06_, S07, S07_, S08, S08_, S09, S10, S11, S11_, S12, S12_,
  SHIFT, SHIFT_, SR_, WGA_
);
defparam iA12.GATE_DELAY = GATE_DELAY;

A13 iA13 (
  rst, ALTEST, ALTM, BMAGZM, CCH33, CDUXD, CDUYD, CDUZD, CGA13, CON2, CTROR,
  CT_, DLKRPT, DRPRST, EMSD, ERRST, F05A_, F05B_, F07A, F07B_, F08B, F10A_,
  F10B, F14B, F14H, FLTOUT, FS01, FS10, G01A, G01A_, G16A_, GOJAM, GYROD,
  IIP, IIP_, INKL, INLNKM, INLNKP, MSTRT, NHALGA, NHVFAL, NOTEST, OTLNKM,
  P02, P02_, P03, P03_, PALE, PIPAFL, RNRADM, RNRADP, SB0_, SB2_, SBY, SCAFAL,
  SHAFTD, STNDBY_, STRT2, SUMA16_, SUMB16_, T03_, T04_, T09_, T10, T10_,
  TC0, TCF0, TEMPIN_, THRSTD, TMPOUT, TRUND, VFAIL, WATCHP, XT0, XT1, d2FSFAL,
  CON3, CTPLS_, DOFILT, FILTIN, MCTRAL_, MOSCAL_, MPIPAL_, MRPTAL_, MSCAFL_,
  MTCAL_, MVFAIL_, MWARNF_, SCADBL, WARN, XT0_, XT1_, AGCWAR, ALGA, CGCWAR,
  CKTAL_, DLKPLS, F08B_, G16SW_, MSTRTP, OSCALM, RESTRT, SBYEXT, STRT1, SYNC14_,
  SYNC4_, TMPCAU
);
defparam iA13.GATE_DELAY = GATE_DELAY;

A14 iA14 (
  rst, BR12B, CGA14, CHINC, CLEARA, CLEARB, CLEARC, CLEARD, DV3764, GOJ1,
  GOJAM, INOUT, MAMU, MNHSBF, MP1, NISQL_, PHS2_, PHS3_, PHS4_, PSEUDO, R1C_,
  RB1_, RSC_, RT_, S01, S01_, S02, S02_, S03, S03_, S04, S04_, S05, S05_,
  S06, S06_, S07, S07_, S08, S08_, S09, S09_, S11, S12, SBY, SCAD, SCAD_,
  STRT2, T01, T01_, T02_, T03, T03_, T04_, T05, T05_, T06, T06_, T07, T07_,
  T08, T08_, T09, T10, T10_, T11, T12A, T12_, TCSAJ3, TIMR, WHOMP_, WL11,
  WL16, WSC_, BR12B_, CLROPE, ERAS, IHENV, ILP, ILP_, NOTEST_, RESETA, RESETB,
  RESETC, RESETD, REX, REY, RILP1, RILP1_, SBE, SBF, SBYREL_, SETAB, SETCD,
  SETEK, WEX, WEY, WL11_, WL16_, XB0, XB0E, XB1, XB1E, XB2E, XB3, XB3E, XB4E,
  XB5, XB5E, XB6, XB6E, XB7E, XT0E, XT1E, XT2E, XT3E, XT4E, XT5E, XT6E, XT7E,
  YB0E, YB1E, YB2E, YB3E, ZID, CXB1_, ERAS_, FNERAS_, NOTEST, R1C, RB1, REDRST,
  ROP_, RSCG_, RSTK_, SBESET, SBFSET, SETAB_, SETCD_, STBE, STBF, STRGAT,
  TPARG_, TPGE, TPGF, WHOMPA, WSCG_, XB0_, XB1_, XB2, XB2_, XB3_, XB4, XB4_,
  XB5_, XB6_, XB7, XB7_, XT0, XT0_, XT1, XT1_, XT2, XT2_, XT3, XT3_, XT4,
  XT4_, XT5, XT5_, XT6, XT6_, XT7, XT7_, YB0, YB0_, YB1, YB1_, YB2, YB2_,
  YB3, YB3_
);
defparam iA14.GATE_DELAY = GATE_DELAY;

A15 iA15 (
  rst, C32M, C32P, C33M, C33P, C34M, C34P, C35M, C35P, C36M, C36P, C37M,
  C40M, C41M, C42M, C43M, C44M, CA2_, CA3_, CAD1, CAD2, CAD3, CEBG, CFBG,
  CGA15, DLKPLS, E5, E6, E7_, GOJAM, HNDRPT, INCSET_, KRPT, KYRPT1, KYRPT2,
  MKRPT, OVF_, R6, RADRPT, RB1F, RBBEG_, REBG_, RFBG_, RRPA, RSTRT, S10,
  S10_, S11_, S12_, STRGAT, SUMA01_, SUMA02_, SUMA03_, SUMA11_, SUMA12_,
  SUMA13_, SUMA14_, SUMA16_, SUMB01_, SUMB02_, SUMB03_, SUMB11_, SUMB12_,
  SUMB13_, SUMB14_, SUMB16_, T10, T12A, U2BBKG_, UPRUPT, WBBEG_, WEBG_, WFBG_,
  WL01_, WL02_, WL03_, WL09_, WL10_, WL11_, WL12_, WL13_, WL14_, WL16_, WOVR,
  XB0_, XB1_, XB4_, XB6_, XB7_, XT0_, XT1_, XT2_, XT3_, XT4_, XT5_, ZOUT_,
  BBK1, BBK2, BBK3, DNRPTA, F11, F11_, F12, F12_, F13, F13_, F14, F14_, F15,
  F15_, F16, F16_, HIMOD, KRPTA_, LOMOD, PRPOR1, PRPOR2, PRPOR3, PRPOR4,
  RL01_, RL02_, RL03_, RL09_, RL10_, RL11_, RL12_, RL13_, RL14_, RL16_, ROPER,
  ROPES, ROPET, RPTA12, RPTAD3, RRPA1_, STR14, STR19, STR210, STR311, STR412,
  STR58, STR912, BK16, DRPRST, EB10, EB10_, EB11, EB11_, EB9, EB9_, FB11,
  FB11_, FB12, FB12_, FB13, FB13_, FB14, FB14_, FB16, FB16_, KY1RST, KY2RST,
  MCDU, MCDU_, MINC, MINC_, PCDU, PCDU_, RPTAD4, RPTAD5, RPTAD6, RUPTOR_,
  T6RPT, WOVR_
);
defparam iA15.GATE_DELAY = GATE_DELAY;

A16 iA16 (
  rst, CCH11, CCHG_, CGA16, CH0705, CH0706, CH0707, CH1501, CH1502, CH1503,
  CH1504, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207, CH3208,
  CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_, CHWL08_,
  CHWL09_, CHWL10_, CHWL11_, CHWL12_, CHWL13_, CHWL14_, FLASH, FLASH_, GOJAM,
  RCH11_, WCH11_, WCHG_, XB2_, XB5_, XB6_, XT0_, XT1_, CCH12, CH1207, CHOR01_,
  CHOR02_, CHOR03_, CHOR04_, CHOR05_, CHOR06_, CHOR07_, CHOR08_, RCH12_,
  WCH12_, CCH05, CCH06, CH1208, CH1209, CH1210, CH1211, CH1212, CH1213, CH1214,
  COARSE, COMACT, DISDAC, ENERIM, ENEROP, ISSWAR, KYRLS, MROLGT, OPEROR,
  OT1207, OT1207_, RCH05_, RCH06_, RCmXmP, RCmXmY, RCmXpP, RCmXpY, RCmYmR,
  RCmYpR, RCmZmR, RCmZpR, RCpXmP, RCpXmY, RCpXpP, RCpXpY, RCpYmR, RCpYpR,
  RCpZmR, RCpZpR, S4BOFF, S4BSEQ, S4BTAK, STARON, TMPOUT, TVCNAB, UPLACT,
  VNFLSH, WCH05_, WCH06_, ZEROPT, ZIMCDU, ZOPCDU
);
defparam iA16.GATE_DELAY = GATE_DELAY;

A17 iA17 (
  rst, AGCWAR, CCHG_, CDUFAL, CGA17, CH1113, CH1213, CH1214, CH1301, CH1302,
  CH1303, CH1304, CH1305, CH1306, CH1307, CH1308, CH1309, CH1310, CH1311,
  CH1316, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406, CH1407, CH1408,
  CH1409, CH1410, CH1411, CH1412, CH1413, CH1414, CH1416, CH3310, CH3312,
  CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_, CHWL08_,
  CHWL09_, CHWL10_, CHWL11_, CHWL12_, CHWL13_, CHWL14_, CHWL16_, CTLSAT,
  F05A_, F05B_, F05D, FREFUN, GCAPCL, GOJAM, GUIREL, HOLFUN, IMUCAG, IMUFAL,
  IMUOPR, IN3008, IN3212, IN3213, IN3214, IN3216, IN3301, ISSTOR, LEMATT,
  LFTOFF, LRRLSC, LVDAGD, MANRmP, MANRmR, MANRmY, MANRpP, MANRpR, MANRpY,
  MNIMmP, MNIMmR, MNIMmY, MNIMpP, MNIMpR, MNIMpY, OPCDFL, OPMSW2, OPMSW3,
  OSCALM, PCHGOF, PIPAFL, ROLGOF, RRPONA, RRRLSC, S01, S02, S4BSAB, SMSEPR,
  SPSRDY, STRPRS, TEMPIN, TPOR_, TRANmX, TRANmY, TRANmZ, TRANpX, TRANpY,
  TRANpZ, TRST10, TRST9, ULLTHR, WCH13_, WCHG_, XB0_, XB1_, XB2_, XB3_, XT1_,
  XT3_, ZEROP, CHOR01_, CHOR02_, CHOR03_, CHOR04_, CHOR05_, CHOR06_, CHOR07_,
  CHOR08_, CHOR09_, CHOR10_, CHOR11_, CHOR12_, CHOR13_, CHOR14_, CHOR16_,
  RCH33_, XB0, CCH10, CCH11, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206,
  CH3207, CH3208, CH3209, CH3210, CH3313, CH3314, CH3316, HNDRPT, RCH10_,
  RCH11_, RCH30_, RCH31_, RCH32_, RLYB01, RLYB02, RLYB03, RLYB04, RLYB05,
  RLYB06, RLYB07, RLYB08, RLYB09, RLYB10, RLYB11, RYWD12, RYWD13, RYWD14,
  RYWD16, TRP31A, TRP31B, TRP32, WCH10_, WCH11_
);
defparam iA17.GATE_DELAY = GATE_DELAY;

A18 iA18 (
  rst, ALTEST, CAURST, CCH13, CCH33, CGA18, CH1111, CH1112, CH1114, CH1116,
  CH1211, CH1212, CH1216, CH3311, CH3313, CH3314, CH3316, CHAT11, CHAT12,
  CHAT13, CHAT14, CHBT11, CHBT12, CHBT13, CHBT14, CHOR11_, CHOR12_, CHOR13_,
  CHOR16_, CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL11_, DKEND, F09A_, F09B,
  F09B_, F09D, F10A, F10A_, F17A, F17B, F5ASB2_, F5BSB2_, GOJAM, GTRST_,
  GTSET_, LRIN0, LRIN1, MAINRS, MARK, MKEY1, MKEY2, MKEY3, MKEY4, MKEY5,
  MRKREJ, MRKRST, NAVRST, NKEY1, NKEY2, NKEY3, NKEY4, NKEY5, RCH13_, RCH33_,
  RCHG_, RRIN0, RRIN1, SB0_, SB2_, SBYBUT, STOP, T05, T11, TEMPIN, W1110,
  WCH13_, XB5_, XB6_, XT1_, CHOR14_, F17A_, F17B_, HERB, TPORA_, TPOR_, CH11,
  CH12, CH13, CH1301, CH1302, CH1303, CH1304, CH1311, CH14, CH1501, CH1502,
  CH1503, CH1504, CH1505, CH16, CH1601, CH1602, CH1603, CH1604, CH1605, CH1606,
  CH1607, CH3312, CNTOF9, DLKRPT, END, ERRST, F10AS0, KYRPT1, KYRPT2, LRRANG,
  LRSYNC, LRXVEL, LRYVEL, LRZVEL, MKRPT, RADRPT, RCH15_, RCH16_, RNRADM,
  RNRADP, RRRANG, RRRARA, RRSYNC, SBY, SBYLIT, STNDBY, STNDBY_, TEMPIN_
);
defparam iA18.GATE_DELAY = GATE_DELAY;

A19 iA19 (
  rst, BLKUPL_, BMGXM, BMGXP, BMGYM, BMGYP, BMGZM, BMGZP, BR1, BR1_, C45R,
  CA2_, CA4_, CA5_, CA6_, CCH11, CCH13, CCH14, CCHG_, CGA19, CHWL01_, CHWL02_,
  CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_, CHWL08_, CHWL09_, CHWL10_,
  CHWL11_, CHWL12_, CNTRSB_, CSG, CXB0_, CXB7_, F04A, F05A_, F05B_, F06B,
  F07B, F07C_, F07D_, F09B, F10A, F10B, F7CSB1_, FS10, GATEX_, GATEY_, GATEZ_,
  GOJAM, GTONE, GTSET, GTSET_, MOUT_, OVF_, POUT_, RCH11_, RCH13_, RCH14_,
  RCH33_, SB0_, SB1_, SB2_, SHINC_, SIGNX, SIGNY, SIGNZ, T06_, T6ON_, UPL0,
  UPL1, WCH11_, WCH13_, WCH14_, WOVR_, XB3_, XB5_, XB6_, XB7_, XLNK0, XLNK1,
  XT3_, ZOUT_, BLKUPL, C45R_, F5ASB0_, F5ASB2, F5ASB2_, UPL0_, UPL1_, XLNK0_,
  XLNK1_, ALRT0, ALRT1, ALT0, ALT1, ALTM, ALTSNC, BMAGXM, BMAGXP, BMAGYM,
  BMAGYP, BMAGZM, BMAGZP, CCH33, CH1109, CH1110, CH1111, CH1112, CH1305,
  CH1306, CH1308, CH1309, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406,
  CH1407, CH1408, CH1409, CH1410, CH3310, CH3311, EMSD, EMSm, EMSp, F06B_,
  F09B_, F10A_, F10B_, F5ASB0, F5BSB2, F5BSB2_, FF1109, FF1109_, FF1110,
  FF1110_, FF1111, FF1111_, FF1112, FF1112_, GYENAB, GYROD, GYRRST, GYRSET,
  GYXM, GYXP, GYYM, GYYP, GYZM, GYZP, INLNKM, INLNKP, OTLNK0, OTLNK1, OTLNKM,
  RHCGO, SH3MS_, T1P, T2P, T3P, T4P, T5P, T6P, THRSTD, THRSTm, THRSTp, UPRUPT,
  W1110
);
defparam iA19.GATE_DELAY = GATE_DELAY;

A20 iA20 (
  rst, BKTF_, CA5_, CDUXD, CDUXM, CDUXP, CDUYD, CDUYM, CDUYP, CDUZD, CDUZM,
  CDUZP, CG26, CGA20, CXB0_, CXB1_, CXB5_, CXB6_, OCTAD2, OCTAD3, OCTAD4,
  OCTAD6, PIPXM, PIPXP, PIPYM, PIPYP, PIPZM, PIPZP, RSSB, SHAFTD, SHAFTM,
  SHAFTP, T1P, T2P, T3P, T4P, T5P, T6P, THRSTD, TRNM, TRNP, TRUND, XB2, XB3,
  XB4, XB7, CA2_, CA3_, CA4_, CG11, CG12, CG14, CG21, CG22, CG24, CXB2_,
  CXB3_, CXB4_, CXB7_, C24A, C24R, C25A, C25R, C26A, C26R, C27A, C27R, C30A,
  C30R, C31A, C31R, C32A, C32M, C32P, C32R, C33A, C33M, C33P, C33R, C34A,
  C34M, C34P, C34R, C35A, C35M, C35P, C35R, C36A, C36M, C36P, C36R, C37A,
  C37M, C37P, C37R, C40A, C40M, C40P, C40R, C41A, C41M, C41P, C41R, C50A,
  C50R, C51A, C51R, C52A, C52R, C53A, C53R, C54A, C54R, C55A, C55R, CA6_,
  CG13, CG23
);
defparam iA20.GATE_DELAY = GATE_DELAY;

A21 iA21 (
  rst, ALTM, BMAGXM, BMAGXP, BMAGYM, BMAGYP, BMAGZM, BMAGZP, C24A, C25A,
  C26A, C27A, C30A, C31A, C32A, C33A, C34A, C35A, C36A, C37A, C40A, C41A,
  C50A, C51A, C52A, C53A, C54A, C55A, CA6_, CG13, CG23, CGA21, CT, CXB2_,
  CXB3_, CXB4_, CXB7_, DOSCAL, EMSD, FS17, GNHNC, GOJAM, GYROD, INLNKM, INLNKP,
  MLDCH, MLOAD, MNHNC, MRDCH, MREAD, NISQL_, OCTAD4, OCTAD5, OTLNKM, PHS2_,
  PHS3_, PHS4_, PSEUDO, RNRADM, RNRADP, RQ, RSCT_, ST0_, ST1_, STD2, T02_,
  T07_, T10_, T11_, T12A, T12_, XB0, XB5, XB6, BKTF_, C42A, C43A, C44A, C45A,
  C45M, C45P, C46A, C46M, C46P, C47A, C56A, C57A, C60A, CA4_, CA5_, CG15,
  CG16, CHINC, CHINC_, CTROR_, CXB0_, CXB5_, CXB6_, DINC, INCSET_, INKBT1,
  INOTLD, INOTRD, MINKL, MREQIN, RSSB, SCAS17, d32004K, C42M, C42P, C42R,
  C43M, C43P, C43R, C44M, C44P, C44R, C45R, C46R, C47R, C56R, C57R, C60R,
  CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CG26, CTROR, DINCNC_, DINC_, FETCH0,
  FETCH0_, FETCH1, INKL, INKL_, MON_, MONpCH, RQ_, SHANC, SHANC_, SHINC,
  SHINC_, STFET1_, STORE1, STORE1_, d30SUM, d50SUM
);
defparam iA21.GATE_DELAY = GATE_DELAY;

A22 iA22 (
  rst, CCH34, CCH35, CCHG_, CGA22, CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL05_,
  CHWL06_, CHWL07_, CHWL08_, CHWL09_, CHWL10_, CHWL11_, CHWL12_, CHWL13_,
  CHWL14_, CHWL16_, DKBSNC, DKSTRT, END, F12B, FS13, FS14, GOJAM, HIGH0_,
  HIGH1_, HIGH2_, HIGH3_, PC15_, WCH34_, WCH35_, WCHG_, XB3_, XB4_, XT1_,
  BSYNC_, CCH13, DATA_, DKCTR2, DKCTR3, DKCTR3_, DKDAT_, DLKCLR, F12B_, FS13_,
  LOW0_, LOW1_, LOW2_, LOW3_, LOW4_, LOW5_, LOW6_, LOW7_, ORDRBT, RCH13_,
  RDOUT_, WCH13_, WDORDR, WRD1B1, WRD1BP, WRD2B2, WRD2B3, ADVCTR, CCH14,
  CH1307, DKCTR1, DKCTR1_, DKCTR2_, DKCTR4, DKCTR4_, DKCTR5, DKCTR5_, DKDATA,
  DKDATB, F14H, RCH14_, WCH14_, d16CNT, d1CNT, d32CNT
);
defparam iA22.GATE_DELAY = GATE_DELAY;

A23 iA23 (
  rst, BOTHZ, CCH11, CCH12, CCH13, CCH14, CCH33, CCHG_, CGA23, CH1109, CH1110,
  CH1208, CH1209, CH1210, CH1505, CH1601, CH1602, CH1603, CH1604, CH1605,
  CH1606, CH1607, CH3209, CH3210, CHAT01, CHAT02, CHAT03, CHAT04, CHAT05,
  CHAT06, CHAT07, CHAT08, CHAT09, CHAT10, CHBT01, CHBT02, CHBT03, CHBT04,
  CHBT05, CHBT06, CHBT07, CHBT08, CHBT09, CHBT10, CHOR01_, CHOR02_, CHOR03_,
  CHOR04_, CHOR05_, CHOR06_, CHOR07_, CHOR08_, CHOR09_, CHOR10_, CHWL01_,
  CHWL05_, CHWL06_, CHWL07_, CHWL08_, CHWL10_, CHWL11_, CHWL12_, CHWL13_,
  CHWL14_, CHWL16_, F18AX, F18B, F5ASB0_, F5ASB2, F5ASB2_, FUTEXT, GOJAM,
  HIGH3_, LOW6_, LOW7_, MISSZ, MOUT, NOZM, NOZP, OCTAD5, PC15_, PHS4_, PIPGXm,
  PIPGXp, PIPGYm, PIPGYp, POUT, RCH11_, RCH12_, RCH13_, RCH14_, RCHG_, T07_,
  T6RPT, WCH11_, WCH12_, WCH13_, WCH14_, WCHG_, XB0_, XB1_, XB2_, XB3_, XB4_,
  XB5_, XB7_, XT0_, XT3_, ZOUT, BOTHX, BOTHY, CH1108, DATA_, F18B_, MISSX,
  MISSY, MOUT_, NOXM, NOXP, NOYM, NOYP, POUT_, T7PHS4, ZOUT_, ALTEST, CCH07,
  CCH34, CCH35, CDUXD, CDUXDM, CDUXDP, CDUYD, CDUYDM, CDUYDP, CDUZD, CDUZDM,
  CDUZDP, CH01, CH02, CH03, CH04, CH05, CH06, CH07, CH0705, CH0706, CH0707,
  CH08, CH09, CH10, CH1113, CH1114, CH1116, CH1216, CH1310, CH1316, CH1411,
  CH1412, CH1413, CH1414, CH1416, E5, E6, E7_, ISSTDC, OT1108, OT1113, OT1114,
  OT1116, PIPAFL, PIPXM, PIPXP, PIPYM, PIPYP, RCH07_, SHAFTD, SHFTDM, SHFTDP,
  T6ON_, T7PHS4_, TRNDM, TRNDP, TRUND, WCH07_, WCH34_, WCH35_
);
defparam iA23.GATE_DELAY = GATE_DELAY;

A24 iA24 (
  rst, A15_, A16_, BMAGXM, BMAGXP, BMAGYM, BMAGYP, BMAGZP, CA6_, CDUXM, CDUXP,
  CDUYM, CDUYP, CDUZM, CDUZP, CGA24, CI_, CT, CT_, DKCTR4, DKCTR4_, DKCTR5,
  DKCTR5_, F01A, F01B, F02B, F03B_, F04B, F05A, F05B, F06B_, F07A_, F07B,
  F08B_, F09A, F17A, F17B, F18AX, F5ASB0, F5ASB2, FF1109_, FF1110_, FF1111_,
  FF1112_, FS02, FS03, FS04, FS05, FS06, FS06_, FS07A, FS07_, FS08, FS08_,
  FS09, FS16, FS17, GOJAM_, IC11, MP3, NISQ_, OCTAD2, OCTAD3, ODDSET_, PIPGZm,
  PIPGZp, PIPXM, PIPXP, PIPYM, PIPYP, RCH_, RSCT, RT_, RUSG_, SB0, SB1, SB2,
  SB4, SHAFTM, SHAFTP, SUMA15_, SUMB15_, T01DC_, T02, T06, T08, T09DC_, T1P,
  T2P, T3P, T4P, T5P, T6P, TRNM, TRNP, U2BBK, WCH_, WL01, WL02, WL03, WL04,
  WL05, WL06, WL07, WL08, WL09, WL10, WL11, WL12, WL13, WL14, WL16, WT_,
  XB3_, XB4_, XB7_, XT0_, CA2_, CA3_, CTPLS_, F05A_, F05B_, F07B_, F5ASB0_,
  F5ASB2_, FS05_, GOJAM, MNISQ, MON800, MRCH, MWATCH_, MWCH, OUTCOM, PIPZM,
  PIPZP, SB0_, SB1_, SB2_, T01, T02_, T09, BOTHZ, CCHG_, CDUCLK, CDUSTB_,
  CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_, CHWL08_,
  CHWL09_, CHWL10_, CHWL11_, CHWL12_, CHWL13_, CHWL14_, CHWL16_, CI, CNTRSB_,
  ELSNCM, ELSNCN, F04B_, F05D, F07C_, F07D_, F09A_, F09D, F7CSB1_, FLASH,
  FLASH_, FS09_, GTONE, GTRST, GTSET, GTSET_, HIGH0_, HIGH1_, HIGH2_, HIGH3_,
  IC11_, LRRST, MISSZ, NISQ, NOZM, NOZP, ONE, OT1110, OT1111, OT1112, OVNHRP,
  PHS3_, PIPASW, PIPDAT, PIPINT, PIPPLS_, RCHAT_, RCHBT_, RCHG_, RRRST, RSCT_,
  U2BBKG_, US2SG, WATCH, WATCHP, WATCH_, WCHG_, d12KPPS, d25KPPS, d3200A,
  d3200B, d3200C, d3200D, d800RST, d800SET
);
defparam iA24.GATE_DELAY = GATE_DELAY;

A99 iA99 (
  rst, GEM01, GEM02, GEM03, GEM04, GEM05, GEM06, GEM07, GEM08, GEM09, GEM10,
  GEM11, GEM12, GEM13, GEM14, GEM16, GEMP, IL01, IL02, IL03, IL04, IL05,
  IL06, IL07, RESETD, REX, REY, RSTKX_, RSTKY_, SBE, SBF, SETAB, SETCD, SETEK,
  STR412, WEX, WEY, XB1E, XB2E, XB4E, XB6E, XT1E, XT2E, XT4E, XT5E, YB1E,
  YB2E, YT1E, YT2E, YT4E, CLROPE, HIMOD, LOMOD, RESETA, RESETB, RESETC, ROPER,
  ROPES, ROPET, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08, SA09, SA10,
  SA11, SA12, SA13, SA14, SA16, SAP, STR14, STR19, STR210, STR311, STR58,
  STR912, XB3E, XB5E, XB7E, XT3E, XT6E, XT7E, YB3E, YT3E, YT5E, YT6E, YT7E,
  ZID
);
defparam iA99.GATE_DELAY = GATE_DELAY;

A52 iA52 (
  rst, p4SW, MCTRAL_, MPAL_, MRCH, MRPTAL_, MSCAFL_, MSCDBL_, MT01, MT05,
  MT12, MTCAL_, MVFAIL_, MWATCH_, MWCH, MWL01, MWL02, MWL03, MWL04, MWL05,
  MWL06, MWSG, DBLTST, DOSCAL, MAMU, MDT01, MDT02, MDT03, MDT04, MDT05, MDT06,
  MDT07, MDT08, MDT09, MDT10, MDT11, MDT12, MDT13, MDT14, MDT15, MDT16, MLDCH,
  MLOAD, MNHNC, MNHRPT, MNHSBF, MONPAR, MONWBK, MRDCH, MREAD, MSBSTP, MSTP,
  MSTRT, MTCSAI, NHALGA
);
defparam iA52.GATE_DELAY = GATE_DELAY;

endmodule
