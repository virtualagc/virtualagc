`timescale 1ns/1ps
`default_nettype none

module memory_timing_addressing(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, STRT2, PHS2_n, PHS3_n, PHS4_n, T01, T01_n, T02_n, T03, T03_n, T04_n, T05, T05_n, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T12_n, T12A, S01, S01_n, S02, S02_n, S03, S03_n, S04, S04_n, S05, S05_n, S06, S06_n, S07, S07_n, S08, S08_n, S09, S09_n, S10_n, S11, S12, EB9, EB10, EB11_n, CHINC, DV3764, GOJ1, INOUT, MP1, TCSAJ3, SCAD, TIMR, MAMU, MNHSBF, STBE, STBF, SBF, STRGAT, TPARG_n, XB0, XB0_n, XB1, XB1_n, XB2, XB2_n, XB3, XB3_n, XB4, XB4_n, XB5, XB5_n, XB6, XB6_n, XB7, XB7_n, XT0_n, XT1_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n, SETAB, SETCD, RESETA, RESETB, RESETC, RESETD, CLROPE, IL01, IL02, IL03, IL04, IL05, IL06, IL07, SBE, SETEK, RSTKX_n, RSTKY_n, REX, REY, WEX, WEY, ZID, XB7E, XB1E, XB2E, XB3E, XB4E, XB5E, XB6E, XT7E, XT1E, XT2E, XT3E, XT4E, XT5E, XT6E, YB3E, YB1E, YB2E, YT7E, YT1E, YT2E, YT3E, YT4E, YT5E, YT6E);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire CHINC;
    output wire CLROPE;
    input wire DV3764;
    input wire EB10;
    input wire EB11_n;
    input wire EB9;
    input wire GOJ1;
    input wire GOJAM;
    output wire IL01;
    output wire IL02;
    output wire IL03;
    output wire IL04;
    output wire IL05;
    output wire IL06;
    output wire IL07;
    input wire INOUT;
    input wire MAMU;
    input wire MNHSBF;
    input wire MP1;
    input wire PHS2_n;
    input wire PHS3_n;
    input wire PHS4_n;
    output wire RESETA;
    output wire RESETB;
    output wire RESETC;
    output wire RESETD;
    output wire REX;
    output wire REY;
    output wire RSTKX_n;
    output wire RSTKY_n;
    input wire S01;
    input wire S01_n;
    input wire S02;
    input wire S02_n;
    input wire S03;
    input wire S03_n;
    input wire S04;
    input wire S04_n;
    input wire S05;
    input wire S05_n;
    input wire S06;
    input wire S06_n;
    input wire S07;
    input wire S07_n;
    input wire S08;
    input wire S08_n;
    input wire S09;
    input wire S09_n;
    input wire S10_n;
    input wire S11;
    input wire S12;
    output wire SBE;
    output wire SBF;
    input wire SCAD;
    output wire SETAB;
    output wire SETCD;
    output wire SETEK;
    output wire STBE;
    output wire STBF;
    output wire STRGAT;
    input wire STRT2;
    input wire T01;
    input wire T01_n;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04_n;
    input wire T05;
    input wire T05_n;
    input wire T06;
    input wire T06_n;
    input wire T07;
    input wire T07_n;
    input wire T08;
    input wire T08_n;
    input wire T09;
    input wire T10;
    input wire T10_n;
    input wire T11;
    input wire T12A;
    input wire T12_n;
    input wire TCSAJ3;
    input wire TIMR;
    output wire TPARG_n;
    output wire WEX;
    output wire WEY;
    output wire XB0;
    output wire XB0_n;
    output wire XB1;
    output wire XB1E;
    output wire XB1_n;
    output wire XB2;
    output wire XB2E;
    output wire XB2_n;
    output wire XB3;
    output wire XB3E;
    output wire XB3_n;
    output wire XB4;
    output wire XB4E;
    output wire XB4_n;
    output wire XB5;
    output wire XB5E;
    output wire XB5_n;
    output wire XB6;
    output wire XB6E;
    output wire XB6_n;
    output wire XB7;
    output wire XB7E;
    output wire XB7_n;
    output wire XT0_n;
    output wire XT1E;
    output wire XT1_n;
    output wire XT2E;
    output wire XT2_n;
    output wire XT3E;
    output wire XT3_n;
    output wire XT4E;
    output wire XT4_n;
    output wire XT5E;
    output wire XT5_n;
    output wire XT6E;
    output wire XT6_n;
    output wire XT7E;
    output wire YB0_n;
    output wire YB1E;
    output wire YB2E;
    output wire YB3E;
    output wire YT0_n;
    output wire YT1E;
    output wire YT2E;
    output wire YT3E;
    output wire YT4E;
    output wire YT5E;
    output wire YT6E;
    output wire YT7E;
    output wire ZID;
    wire __A14_1__CLEARA;
    wire __A14_1__CLEARB;
    wire __A14_1__CLEARC;
    wire __A14_1__CLEARD;
    wire __A14_1__ERAS; //FPGA#wand
    wire __A14_1__ERAS_n;
    wire __A14_1__FNERAS_n;
    wire __A14_1__IHENV;
    wire __A14_1__REDRST;
    wire __A14_1__ROP_n;
    wire __A14_1__RSTK_n;
    wire __A14_1__S08A;
    wire __A14_1__S08A_n;
    wire __A14_1__SBESET;
    wire __A14_1__SBFSET; //FPGA#wand
    wire __A14_1__SETAB_n;
    wire __A14_1__SETCD_n;
    wire __A14_1__TPGE; //FPGA#wand
    wire __A14_1__TPGF; //FPGA#wand
    wire __A14_2__EAD09;
    wire __A14_2__EAD09_n;
    wire __A14_2__EAD10;
    wire __A14_2__EAD10_n;
    wire __A14_2__EAD11;
    wire __A14_2__EAD11_n;
    wire __A14_2__IL01_n;
    wire __A14_2__IL02_n;
    wire __A14_2__IL03_n;
    wire __A14_2__IL04_n;
    wire __A14_2__IL05_n;
    wire __A14_2__IL06_n;
    wire __A14_2__IL07_n;
    wire __A14_2__ILP;
    wire __A14_2__ILP_n;
    wire __A14_2__RILP1;
    wire __A14_2__RILP1_n;
    wire __A14_2__XB0E;
    wire __A14_2__XT0;
    wire __A14_2__XT0E;
    wire __A14_2__XT1;
    wire __A14_2__XT2;
    wire __A14_2__XT3;
    wire __A14_2__XT4;
    wire __A14_2__XT5;
    wire __A14_2__XT6;
    wire __A14_2__XT7;
    wire __A14_2__XT7_n;
    wire __A14_2__YB0;
    wire __A14_2__YB0E;
    wire __A14_2__YB1;
    wire __A14_2__YB1_n;
    wire __A14_2__YB2;
    wire __A14_2__YB2_n;
    wire __A14_2__YB3;
    wire __A14_2__YB3_n;
    wire __A14_2__YT0;
    wire __A14_2__YT0E;
    wire __A14_2__YT1;
    wire __A14_2__YT1_n;
    wire __A14_2__YT2;
    wire __A14_2__YT2_n;
    wire __A14_2__YT3;
    wire __A14_2__YT3_n;
    wire __A14_2__YT4;
    wire __A14_2__YT4_n;
    wire __A14_2__YT5;
    wire __A14_2__YT5_n;
    wire __A14_2__YT6;
    wire __A14_2__YT6_n;
    wire __A14_2__YT7;
    wire __A14_2__YT7_n;
    wire net_U14001_Pad10;
    wire net_U14001_Pad11;
    wire net_U14001_Pad12;
    wire net_U14001_Pad13;
    wire net_U14001_Pad4;
    wire net_U14001_Pad9;
    wire net_U14002_Pad10;
    wire net_U14003_Pad11;
    wire net_U14003_Pad5;
    wire net_U14004_Pad12;
    wire net_U14004_Pad13;
    wire net_U14004_Pad6;
    wire net_U14004_Pad8;
    wire net_U14005_Pad12;
    wire net_U14005_Pad13;
    wire net_U14006_Pad6;
    wire net_U14006_Pad8;
    wire net_U14007_Pad1;
    wire net_U14007_Pad10;
    wire net_U14007_Pad12;
    wire net_U14007_Pad13;
    wire net_U14007_Pad4;
    wire net_U14007_Pad9;
    wire net_U14009_Pad10;
    wire net_U14009_Pad11;
    wire net_U14011_Pad10;
    wire net_U14011_Pad13;
    wire net_U14012_Pad11;
    wire net_U14012_Pad4;
    wire net_U14012_Pad9;
    wire net_U14013_Pad12;
    wire net_U14013_Pad6;
    wire net_U14014_Pad11;
    wire net_U14014_Pad13;
    wire net_U14014_Pad5;
    wire net_U14014_Pad9;
    wire net_U14016_Pad12;
    wire net_U14016_Pad13;
    wire net_U14016_Pad6;
    wire net_U14016_Pad8;
    wire net_U14016_Pad9;
    wire net_U14017_Pad1;
    wire net_U14017_Pad12;
    wire net_U14017_Pad13;
    wire net_U14018_Pad10;
    wire net_U14018_Pad11;
    wire net_U14018_Pad12;
    wire net_U14018_Pad3;
    wire net_U14019_Pad11;
    wire net_U14019_Pad6;
    wire net_U14019_Pad8;
    wire net_U14020_Pad13;
    wire net_U14020_Pad3;
    wire net_U14020_Pad6;
    wire net_U14021_Pad1;
    wire net_U14021_Pad12;
    wire net_U14021_Pad2;
    wire net_U14021_Pad6;
    wire net_U14021_Pad8;
    wire net_U14022_Pad10;
    wire net_U14022_Pad13;
    wire net_U14022_Pad4;
    wire net_U14022_Pad8;
    wire net_U14024_Pad12;
    wire net_U14024_Pad13;
    wire net_U14024_Pad3;
    wire net_U14024_Pad6;
    wire net_U14024_Pad8;
    wire net_U14024_Pad9;
    wire net_U14025_Pad10;
    wire net_U14027_Pad11;
    wire net_U14028_Pad5;
    wire net_U14030_Pad10;
    wire net_U14030_Pad13;
    wire net_U14030_Pad2;
    wire net_U14031_Pad4;
    wire net_U14032_Pad12;
    wire net_U14039_Pad13;
    wire net_U14047_Pad4;
    wire net_U14052_Pad12;
    wire net_U14052_Pad13;
    wire net_U14053_Pad11;
    wire net_U14053_Pad8;
    wire net_U14055_Pad11;
    wire net_U14055_Pad2;
    wire net_U14055_Pad5;
    wire net_U14056_Pad12;
    wire net_U14056_Pad6;
    wire net_U14056_Pad8;

    pullup R14001(__A14_1__SBFSET);
    pullup R14002(__A14_1__TPGF);
    pullup R14003(__A14_1__ERAS);
    pullup R14004(__A14_1__TPGE);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14001(__A14_1__ROP_n, S11, S12, net_U14001_Pad4, T08_n, PHS3_n, GND, net_U14001_Pad4, net_U14001_Pad9, net_U14001_Pad10, net_U14001_Pad11, net_U14001_Pad12, net_U14001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14002(net_U14001_Pad10, T09, __A14_1__ROP_n, net_U14001_Pad10, T08, net_U14001_Pad11, GND, net_U14001_Pad12, net_U14001_Pad13, net_U14002_Pad10, TIMR, net_U14001_Pad9, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14003(T01_n, net_U14002_Pad10, net_U14001_Pad13, __A14_1__IHENV, net_U14003_Pad5, __A14_1__SETAB_n, GND, SETAB, __A14_1__SETAB_n, __A14_1__SETCD_n, net_U14003_Pad11, SETCD, __A14_1__SETCD_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14004(TIMR, net_U14002_Pad10, PHS4_n, __A14_1__ROP_n, T10_n, net_U14004_Pad6, GND, net_U14004_Pad8, T05_n, PHS3_n, __A14_1__ROP_n, net_U14004_Pad12, net_U14004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14005(net_U14004_Pad13, net_U14004_Pad12, net_U14004_Pad6, net_U14003_Pad5, S09, net_U14004_Pad13, GND, net_U14004_Pad13, S09_n, net_U14003_Pad11, net_U14004_Pad8, net_U14005_Pad12, net_U14005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14006(net_U14005_Pad13, T08, net_U14005_Pad13, S09, S08, net_U14006_Pad6, GND, net_U14006_Pad8, net_U14005_Pad13, S09, S08_n, net_U14005_Pad12, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14007(net_U14007_Pad1, __A14_1__CLEARA, net_U14006_Pad6, net_U14007_Pad4, __A14_1__CLEARB, net_U14006_Pad8, GND, __A14_1__CLEARC, net_U14007_Pad9, net_U14007_Pad10, __A14_1__CLEARD, net_U14007_Pad12, net_U14007_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14008(net_U14007_Pad1, RESETA, net_U14007_Pad4, RESETB, net_U14007_Pad10, RESETC, GND, RESETD, net_U14007_Pad13, __A14_1__S08A_n, S08, __A14_1__S08A, S08_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14009(net_U14005_Pad13, S08, net_U14005_Pad13, S09_n, S08_n, net_U14007_Pad12, GND, STBF, GOJAM, net_U14009_Pad10, net_U14009_Pad11, net_U14007_Pad9, S09_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14010(__A14_1__CLEARA, __A14_1__SETAB_n, __A14_1__S08A_n, __A14_1__CLEARB, __A14_1__SETAB_n, __A14_1__S08A, GND, __A14_1__SETCD_n, __A14_1__S08A_n, __A14_1__CLEARC, __A14_1__SETCD_n, __A14_1__S08A, __A14_1__CLEARD, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14011(net_U14009_Pad11, STBF, __A14_1__SBFSET, net_U14009_Pad10, T07_n, PHS3_n, GND, T02_n, __A14_1__ROP_n, net_U14011_Pad10, net_U14011_Pad10, STRGAT, net_U14011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14012(net_U14009_Pad11, SBF, __A14_1__ROP_n, net_U14012_Pad4, S07_n, __A14_2__IL07_n, GND, WEX, net_U14012_Pad9, WEY, net_U14012_Pad11, __A14_1__ERAS_n, __A14_1__ERAS, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14013(MNHSBF, MP1, __A14_1__ROP_n, T06_n, DV3764, net_U14013_Pad6, GND, STRGAT, net_U14011_Pad13, T08, GOJAM, net_U14013_Pad12, PHS4_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U14014(net_U14013_Pad12, __A14_1__SBFSET, net_U14013_Pad6, __A14_1__SBFSET, net_U14014_Pad5, __A14_1__TPGF, GND, __A14_1__TPGF, net_U14014_Pad9, __A14_1__ERAS, net_U14014_Pad11, __A14_1__ERAS, net_U14014_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U14015(net_U14014_Pad5, __A14_1__ROP_n, T08_n, DV3764, GOJ1,  , GND,  , GOJAM, TCSAJ3, PHS2_n, MP1, net_U14014_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14016(T02_n, net_U14012_Pad4, net_U14016_Pad13, T03, GOJAM, net_U14016_Pad6, GND, net_U14016_Pad8, net_U14016_Pad9, T07, GOJAM, net_U14016_Pad12, net_U14016_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U14017(net_U14017_Pad1, __A14_1__ROP_n, T10_n, net_U14016_Pad13, net_U14017_Pad1, net_U14016_Pad6, GND, net_U14016_Pad12, net_U14016_Pad8, net_U14016_Pad9, T01, net_U14017_Pad12, net_U14017_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14018(net_U14017_Pad12, net_U14017_Pad13, net_U14018_Pad3, net_U14018_Pad3, T12_n, PHS3_n, GND, T12A, net_U14017_Pad12, net_U14018_Pad10, net_U14018_Pad11, net_U14018_Pad12, net_U14012_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14019(net_U14018_Pad10, TIMR, net_U14018_Pad10, TIMR, net_U14012_Pad11, net_U14019_Pad6, GND, net_U14019_Pad8, TIMR, T11, net_U14019_Pad11, net_U14018_Pad11, net_U14012_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U14020(net_U14012_Pad11, net_U14019_Pad6, net_U14020_Pad3, net_U14019_Pad11, net_U14019_Pad8, net_U14020_Pad6, GND, net_U14019_Pad11, T10, net_U14018_Pad12, T05_n, __A14_1__ERAS_n, net_U14020_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14021(net_U14021_Pad1, net_U14021_Pad2, __A14_1__ERAS_n, PHS3_n, T03_n, net_U14021_Pad6, GND, net_U14021_Pad8, __A14_1__FNERAS_n, T12A, GOJAM, net_U14021_Pad12, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U14022(__A14_1__FNERAS_n, net_U14020_Pad13, net_U14021_Pad8, net_U14022_Pad4, __A14_1__FNERAS_n, T10_n, GND, net_U14022_Pad8, net_U14020_Pad6, net_U14022_Pad10, T02_n, PHS4_n, net_U14022_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14023(T10_n, __A14_1__FNERAS_n, __A14_1__FNERAS_n, T10_n, PHS3_n, net_U14020_Pad6, GND, net_U14022_Pad8, TIMR, net_U14022_Pad13, net_U14022_Pad10, net_U14020_Pad3, PHS4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14024(TIMR, T01, net_U14024_Pad3, GOJAM, __A14_1__REDRST, net_U14024_Pad6, GND, net_U14024_Pad8, net_U14024_Pad9, GOJAM, __A14_1__REDRST, net_U14024_Pad12, net_U14024_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14025(net_U14024_Pad13, net_U14024_Pad12, net_U14022_Pad4, ZID, net_U14024_Pad13, STRT2, GND, __A14_1__ERAS_n, T03_n, net_U14025_Pad10, net_U14025_Pad10, net_U14021_Pad12, net_U14021_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14026(net_U14014_Pad11, TCSAJ3, S11, S12, INOUT,  , GND,  , CHINC, GOJ1, MP1, MAMU, net_U14014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14027(SETEK, STRT2, net_U14021_Pad1, net_U14021_Pad2, T06_n, PHS3_n, GND, net_U14021_Pad6, net_U14024_Pad6, net_U14024_Pad3, net_U14027_Pad11, net_U14024_Pad8, net_U14024_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14028(net_U14024_Pad3, REY, net_U14024_Pad9, REX, net_U14028_Pad5, SBE, GND, __A14_1__RSTK_n, net_U14022_Pad10, RSTKY_n, __A14_1__RSTK_n, RSTKX_n, __A14_1__RSTK_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14029(__A14_1__ERAS_n, T03_n, GOJAM, T05, net_U14028_Pad5, STBE, GND, __A14_1__SBESET, T04_n, __A14_1__ERAS_n, SCAD, net_U14027_Pad11, PHS4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U14030(__A14_1__REDRST, net_U14030_Pad2, T05, net_U14030_Pad2, net_U14030_Pad13, net_U14030_Pad10, GND, net_U14030_Pad2, T06, net_U14030_Pad10, T05_n, PHS3_n, net_U14030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U14031(net_U14028_Pad5, STBE, __A14_1__SBESET, net_U14031_Pad4, T05_n, PHS3_n, GND, __A14_1__TPGF, __A14_1__TPGE, TPARG_n, S07, S08, __A14_2__YB0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14032(SCAD, __A14_1__ERAS_n, S01, S02, S03, XB0, GND, XB1, S01_n, S02, S03, net_U14032_Pad12, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U14033(net_U14032_Pad12, __A14_1__TPGE, net_U14031_Pad4, __A14_1__TPGE,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4
    U74HC04 U14034(XB0, XB0_n, XB0_n, __A14_2__XB0E, XB1, XB1_n, GND, XB1E, XB1_n, XB2_n, XB2, XB2E, XB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14035(S01, S02_n, S01_n, S02_n, S03, XB3, GND, XB4, S01, S02, S03_n, XB2, S03, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14036(XB3, XB3_n, XB3_n, XB3E, XB4, XB4_n, GND, XB4E, XB4_n, XB5_n, XB5, XB5E, XB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14037(S01_n, S02, S01, S02_n, S03_n, XB6, GND, XB7, S01_n, S02_n, S03_n, XB5, S03_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14038(XB6, XB6_n, XB6_n, XB6E, XB7, XB7_n, GND, XB7E, XB7_n, YB0_n, __A14_2__YB0, __A14_2__YB0E, YB0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14039(__A14_2__YB1, S07_n, S08, __A14_2__YB2, S07, S08_n, GND, S07_n, S08_n, __A14_2__YB3, EB9, S10_n, net_U14039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14040(__A14_2__YB1, __A14_2__YB1_n, __A14_2__YB1_n, YB1E, __A14_2__YB2, __A14_2__YB2_n, GND, YB2E, __A14_2__YB2_n, __A14_2__YB3_n, __A14_2__YB3, YB3E, __A14_2__YB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14041(S04, S05, S04_n, S05, S06, __A14_2__XT1, GND, __A14_2__XT2, S04, S05_n, S06, __A14_2__XT0, S06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14042(__A14_2__XT0, XT0_n, XT0_n, __A14_2__XT0E, __A14_2__XT1, XT1_n, GND, XT1E, XT1_n, XT2_n, __A14_2__XT2, XT2E, XT2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14043(S04_n, S05_n, S04, S05, S06_n, __A14_2__XT4, GND, __A14_2__XT5, S04_n, S05, S06_n, __A14_2__XT3, S06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14044(__A14_2__XT3, XT3_n, XT3_n, XT3E, __A14_2__XT4, XT4_n, GND, XT4E, XT4_n, XT5_n, __A14_2__XT5, XT5E, XT5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14045(S04, S05_n, S04_n, S05_n, S06_n, __A14_2__XT7, GND, __A14_2__EAD11, S09_n, S10_n, EB11_n, __A14_2__XT6, S06_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14046(__A14_2__XT6, XT6_n, XT6_n, XT6E, __A14_2__XT7, __A14_2__XT7_n, GND, XT7E, __A14_2__XT7_n, __A14_2__EAD09_n, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14047(__A14_2__EAD09, net_U14039_Pad13, S09_n, net_U14047_Pad4, EB10, S09_n, GND, S10_n, net_U14047_Pad4, __A14_2__EAD10, __A14_2__YB0, __A14_2__YB3, __A14_2__RILP1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14048(__A14_2__EAD11, __A14_2__EAD11_n, __A14_2__YT0, YT0_n, YT0_n, __A14_2__YT0E, GND, __A14_2__YT1_n, __A14_2__YT1, YT1E, __A14_2__YT1_n, __A14_2__YT2_n, __A14_2__YT2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14049(__A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11, __A14_2__YT1, GND, __A14_2__YT2, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD11, __A14_2__YT0, __A14_2__EAD11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14050(__A14_2__YT2_n, YT2E, __A14_2__YT3, __A14_2__YT3_n, __A14_2__YT3_n, YT3E, GND, __A14_2__YT4_n, __A14_2__YT4, YT4E, __A14_2__YT4_n, __A14_2__YT5_n, __A14_2__YT5, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14051(__A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT4, GND, __A14_2__YT5, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT3, __A14_2__EAD11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14052(__A14_2__YT5_n, YT5E, __A14_2__YT6, __A14_2__YT6_n, __A14_2__YT6_n, YT6E, GND, __A14_2__YT7_n, __A14_2__YT7, YT7E, __A14_2__YT7_n, net_U14052_Pad12, net_U14052_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14053(__A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD11_n, __A14_2__YT7, GND, net_U14053_Pad8, net_U14052_Pad13, __A14_2__RILP1, net_U14053_Pad11, __A14_2__YT6, __A14_2__EAD11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14054(net_U14052_Pad13, XB0, XB3, XB5, XB6,  , GND,  , __A14_2__XT0, __A14_2__XT3, __A14_2__XT5, __A14_2__XT6, net_U14053_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14055(net_U14053_Pad11, net_U14055_Pad2, __A14_2__RILP1, __A14_2__RILP1_n, net_U14055_Pad5, net_U14055_Pad11, GND, __A14_2__ILP_n, net_U14055_Pad5, __A14_2__ILP, net_U14055_Pad11, IL01, S01, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14056(net_U14052_Pad12, __A14_2__RILP1, net_U14052_Pad12, __A14_2__RILP1_n, net_U14053_Pad11, net_U14056_Pad6, GND, net_U14056_Pad8, net_U14052_Pad13, __A14_2__RILP1_n, net_U14055_Pad2, net_U14056_Pad12, net_U14055_Pad2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14057(net_U14055_Pad5, net_U14053_Pad8, net_U14056_Pad12, net_U14056_Pad6, net_U14056_Pad8,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14058(S01_n, __A14_2__IL01_n, S02, IL02, S02_n, __A14_2__IL02_n, GND, IL03, S03, __A14_2__IL03_n, S03_n, IL04, S04, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14059(S04_n, __A14_2__IL04_n, S05, IL05, S05_n, __A14_2__IL05_n, GND, IL06, S06, __A14_2__IL06_n, S06_n, IL07, S07, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14060(CLROPE, STRT2, net_U14016_Pad9,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule