// Verilog testbench created by dumbTestbench.py
`timescale 100ns / 1ns

module agc;

reg rst = 1;
reg STRT2 = 1;
initial
  begin
    $dumpfile("agc.lxt2");
    $dumpvars(0, agc);
    # 1 rst = 0;
    # 50 STRT2 = 0;
    # 1000 $finish;
  end

reg CLOCK = 0;
always #2.44140625 CLOCK = !CLOCK;

reg BLKUPL_ = 0, BMGXM = 0, BMGXP = 0, BMGYM = 0, BMGYP = 0, BMGZM = 0,
  BMGZP = 0, BR1 = 0, BR1_ = 0, C45R = 0, CA2_ = 0, CA4_ = 0, CA5_ = 0,
  CA6_ = 0, CCH11 = 0, CCH13 = 0, CCH14 = 0, CCHG_ = 0, CGA19 = 0, CHWL01_ = 0,
  CHWL02_ = 0, CHWL03_ = 0, CHWL04_ = 0, CHWL05_ = 0, CHWL06_ = 0, CHWL07_ = 0,
  CHWL08_ = 0, CHWL09_ = 0, CHWL10_ = 0, CHWL11_ = 0, CHWL12_ = 0, CNTRSB_ = 0,
  CSG = 0, CXB0_ = 0, CXB7_ = 0, F04A = 0, F05A_ = 0, F05B_ = 0, F06B = 0,
  F07B = 0, F07C_ = 0, F07D_ = 0, F09B = 0, F10A = 0, F10B = 0, F7CSB1_ = 0,
  FS10 = 0, GATEX_ = 0, GATEY_ = 0, GATEZ_ = 0, GOJAM = 0, GTONE = 0, GTSET = 0,
  GTSET_ = 0, MOUT_ = 0, OVF_ = 0, POUT_ = 0, RCH11_ = 0, RCH13_ = 0, RCH14_ = 0,
  RCH33_ = 0, SB0_ = 0, SB1_ = 0, SB2_ = 0, SHINC_ = 0, SIGNX = 0, SIGNY = 0,
  SIGNZ = 0, T06_ = 0, T6ON_ = 0, UPL0 = 0, UPL1 = 0, WCH11_ = 0, WCH13_ = 0,
  WCH14_ = 0, WOVR_ = 0, XB3_ = 0, XB5_ = 0, XB6_ = 0, XB7_ = 0, XLNK0 = 0,
  XLNK1 = 0, XT3_ = 0, ZOUT_ = 0;

wire ALRT0, ALRT1, ALT0, ALT1, ALTM, ALTSNC, BLKUPL, BMAGXM, BMAGXP, BMAGYM,
  BMAGYP, BMAGZM, BMAGZP, C45R_, CCH33, CH1109, CH1110, CH1111, CH1112,
  CH1305, CH1306, CH1308, CH1309, CH1401, CH1402, CH1403, CH1404, CH1405,
  CH1406, CH1407, CH1408, CH1409, CH1410, CH3310, CH3311, EMSD, EMSm, EMSp,
  F06B_, F09B_, F10A_, F10B_, F5ASB0, F5ASB0_, F5ASB2, F5ASB2_, F5BSB2,
  F5BSB2_, FF1109, FF1109_, FF1110, FF1110_, FF1111, FF1111_, FF1112, FF1112_,
  GYENAB, GYROD, GYRRST, GYRSET, GYXM, GYXP, GYYM, GYYP, GYZM, GYZP, INLNKM,
  INLNKP, OTLNK0, OTLNK1, OTLNKM, RHCGO, SH3MS_, T1P, T2P, T3P, T4P, T5P,
  T6P, THRSTD, THRSTm, THRSTp, UPL0_, UPL1_, UPRUPT, W1110, XLNK0_, XLNK1_;

A19 iA19 (
  rst, BLKUPL_, BMGXM, BMGXP, BMGYM, BMGYP, BMGZM, BMGZP, BR1, BR1_, C45R,
  CA2_, CA4_, CA5_, CA6_, CCH11, CCH13, CCH14, CCHG_, CGA19, CHWL01_, CHWL02_,
  CHWL03_, CHWL04_, CHWL05_, CHWL06_, CHWL07_, CHWL08_, CHWL09_, CHWL10_,
  CHWL11_, CHWL12_, CNTRSB_, CSG, CXB0_, CXB7_, F04A, F05A_, F05B_, F06B,
  F07B, F07C_, F07D_, F09B, F10A, F10B, F7CSB1_, FS10, GATEX_, GATEY_, GATEZ_,
  GOJAM, GTONE, GTSET, GTSET_, MOUT_, OVF_, POUT_, RCH11_, RCH13_, RCH14_,
  RCH33_, SB0_, SB1_, SB2_, SHINC_, SIGNX, SIGNY, SIGNZ, T06_, T6ON_, UPL0,
  UPL1, WCH11_, WCH13_, WCH14_, WOVR_, XB3_, XB5_, XB6_, XB7_, XLNK0, XLNK1,
  XT3_, ZOUT_, BLKUPL, C45R_, F5ASB0_, F5ASB2, F5ASB2_, UPL0_, UPL1_, XLNK0_,
  XLNK1_, ALRT0, ALRT1, ALT0, ALT1, ALTM, ALTSNC, BMAGXM, BMAGXP, BMAGYM,
  BMAGYP, BMAGZM, BMAGZP, CCH33, CH1109, CH1110, CH1111, CH1112, CH1305,
  CH1306, CH1308, CH1309, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406,
  CH1407, CH1408, CH1409, CH1410, CH3310, CH3311, EMSD, EMSm, EMSp, F06B_,
  F09B_, F10A_, F10B_, F5ASB0, F5BSB2, F5BSB2_, FF1109, FF1109_, FF1110,
  FF1110_, FF1111, FF1111_, FF1112, FF1112_, GYENAB, GYROD, GYRRST, GYRSET,
  GYXM, GYXP, GYYM, GYYP, GYZM, GYZP, INLNKM, INLNKP, OTLNK0, OTLNK1, OTLNKM,
  RHCGO, SH3MS_, T1P, T2P, T3P, T4P, T5P, T6P, THRSTD, THRSTm, THRSTp, UPRUPT,
  W1110
);

initial $timeformat(-9, 0, " ns", 10);
initial $monitor("%t: %d", $time, CLOCK);

endmodule
