`timescale 1ns/1ps
`default_nettype none

module parity_s_register(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, PHS4_n, T02_n, T07_n, T12A, TPARG_n, TSUDO_n, FUTEXT, CGG, CSG, WEDOPG_n, WSG_n, G01, G02, G03, G04, G05, G06, G07, G08, G09, G10, G11, G12, G13, G14, G15, G16, WL01_n, WL02_n, WL03_n, WL04_n, WL05_n, WL06_n, WL07_n, WL08_n, WL09_n, WL10_n, WL11_n, WL12_n, WL13_n, WL14_n, SUMA16_n, SUMB16_n, RAD, SAP, SCAD, OCTAD2, n8XP5, MONPAR, XB0_n, XB1_n, XB2_n, XB3_n, CYL_n, CYR_n, EDOP_n, GINH, SR_n, EXTPLS, INHPLS, RELPLS, G01ED, G02ED, G03ED, G04ED, G05ED, G06ED, G07ED, GEQZRO_n, RADRG, RADRZ, S01, S01_n, S02, S02_n, S03, S03_n, S04, S04_n, S05, S05_n, S06, S06_n, S07, S07_n, S08, S08_n, S09, S09_n, S10, S10_n, S11, S11_n, S12, S12_n, GEMP, G16SW_n, PC15_n, PALE, MGP_n, MSP, MPAL_n);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire CGG;
    input wire CSG;
    output wire CYL_n;
    output wire CYR_n;
    output wire EDOP_n;
    output wire EXTPLS;
    input wire FUTEXT;
    input wire G01;
    output wire G01ED;
    input wire G02;
    output wire G02ED;
    input wire G03;
    output wire G03ED;
    input wire G04;
    output wire G04ED;
    input wire G05;
    output wire G05ED;
    input wire G06;
    output wire G06ED;
    input wire G07;
    output wire G07ED;
    input wire G08;
    input wire G09;
    input wire G10;
    input wire G11;
    input wire G12;
    input wire G13;
    input wire G14;
    input wire G15;
    input wire G16;
    output wire G16SW_n;
    output wire GEMP;
    output wire GEQZRO_n;
    output wire GINH;
    input wire GOJAM;
    inout wire INHPLS; //FPGA#wand
    output wire MGP_n;
    input wire MONPAR;
    output wire MPAL_n; //FPGA#wand
    output wire MSP;
    input wire OCTAD2;
    inout wire PALE; //FPGA#wand
    output wire PC15_n;
    input wire PHS4_n;
    input wire RAD;
    output wire RADRG;
    output wire RADRZ;
    inout wire RELPLS; //FPGA#wand
    output wire S01;
    output wire S01_n;
    output wire S02;
    output wire S02_n;
    output wire S03;
    output wire S03_n;
    output wire S04;
    output wire S04_n;
    output wire S05;
    output wire S05_n;
    output wire S06;
    output wire S06_n;
    output wire S07;
    output wire S07_n;
    output wire S08;
    output wire S08_n;
    output wire S09;
    output wire S09_n;
    output wire S10;
    output wire S10_n;
    output wire S11;
    output wire S11_n;
    output wire S12;
    output wire S12_n;
    input wire SAP;
    input wire SCAD;
    output wire SR_n;
    input wire SUMA16_n;
    input wire SUMB16_n;
    input wire T02_n;
    input wire T07_n;
    input wire T12A;
    input wire TPARG_n;
    input wire TSUDO_n;
    input wire WEDOPG_n;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL07_n;
    input wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WSG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    wire __A12_1__G01A_n;
    wire __A12_1__G16A_n;
    wire __A12_1__GNZRO; //FPGA#wand
    wire __A12_1__PA03;
    wire __A12_1__PA03_n;
    wire __A12_1__PA06;
    wire __A12_1__PA06_n;
    wire __A12_1__PA09;
    wire __A12_1__PA09_n;
    wire __A12_1__PA12;
    wire __A12_1__PA12_n;
    wire __A12_1__PA15;
    wire __A12_1__PA15_n;
    wire __A12_1__PB09;
    wire __A12_1__PB09_n;
    wire __A12_1__PB15;
    wire __A12_1__PB15_n;
    wire __A12_1__PC15;
    wire __A12_1__T7PHS4;
    wire __A12_1__T7PHS4_n;
    wire __A12_1__uG02_n;
    wire __A12_1__uG03_n;
    wire __A12_2__G01A;
    input wire n8XP5;
    wire net_U12001_Pad10;
    wire net_U12001_Pad12;
    wire net_U12002_Pad12;
    wire net_U12002_Pad6;
    wire net_U12002_Pad8;
    wire net_U12003_Pad11;
    wire net_U12003_Pad12;
    wire net_U12003_Pad6;
    wire net_U12003_Pad8;
    wire net_U12004_Pad11;
    wire net_U12004_Pad12;
    wire net_U12005_Pad10;
    wire net_U12005_Pad12;
    wire net_U12005_Pad4;
    wire net_U12005_Pad8;
    wire net_U12006_Pad8;
    wire net_U12007_Pad12;
    wire net_U12007_Pad6;
    wire net_U12007_Pad8;
    wire net_U12008_Pad10;
    wire net_U12008_Pad11;
    wire net_U12008_Pad12;
    wire net_U12008_Pad9;
    wire net_U12009_Pad10;
    wire net_U12009_Pad12;
    wire net_U12009_Pad2;
    wire net_U12009_Pad6;
    wire net_U12009_Pad8;
    wire net_U12011_Pad10;
    wire net_U12011_Pad6;
    wire net_U12011_Pad8;
    wire net_U12012_Pad10;
    wire net_U12012_Pad4;
    wire net_U12013_Pad12;
    wire net_U12013_Pad6;
    wire net_U12013_Pad8;
    wire net_U12014_Pad12;
    wire net_U12014_Pad13;
    wire net_U12015_Pad1;
    wire net_U12015_Pad10;
    wire net_U12015_Pad13;
    wire net_U12015_Pad4;
    wire net_U12016_Pad11;
    wire net_U12016_Pad5;
    wire net_U12017_Pad10;
    wire net_U12017_Pad2;
    wire net_U12017_Pad4;
    wire net_U12017_Pad6;
    wire net_U12017_Pad9;
    wire net_U12019_Pad10;
    wire net_U12019_Pad11;
    wire net_U12019_Pad12;
    wire net_U12019_Pad9;
    wire net_U12020_Pad13;
    wire net_U12022_Pad10;
    wire net_U12022_Pad3;
    wire net_U12022_Pad6;
    wire net_U12022_Pad8;
    wire net_U12023_Pad1;
    wire net_U12023_Pad10;
    wire net_U12023_Pad13;
    wire net_U12025_Pad13;
    wire net_U12026_Pad11;
    wire net_U12026_Pad12;
    wire net_U12026_Pad8;
    wire net_U12028_Pad10;
    wire net_U12028_Pad13;
    wire net_U12028_Pad4;
    wire net_U12029_Pad11;
    wire net_U12029_Pad13;
    wire net_U12029_Pad5;
    wire net_U12029_Pad9;
    wire net_U12030_Pad4;
    wire net_U12031_Pad4;
    wire net_U12032_Pad10;
    wire net_U12032_Pad13;
    wire net_U12032_Pad4;
    wire net_U12033_Pad11;
    wire net_U12033_Pad13;
    wire net_U12033_Pad5;
    wire net_U12033_Pad9;
    wire net_U12034_Pad10;
    wire net_U12034_Pad4;
    wire net_U12035_Pad10;
    wire net_U12036_Pad10;
    wire net_U12036_Pad13;
    wire net_U12036_Pad4;
    wire net_U12037_Pad11;
    wire net_U12037_Pad13;
    wire net_U12037_Pad5;
    wire net_U12037_Pad9;
    wire net_U12038_Pad1;
    wire net_U12038_Pad13;
    wire net_U12039_Pad10;
    wire net_U12039_Pad12;
    wire net_U12039_Pad13;
    wire net_U12040_Pad10;
    wire net_U12040_Pad13;
    wire net_U12040_Pad4;
    wire net_U12041_Pad11;
    wire net_U12041_Pad13;
    wire net_U12042_Pad1;
    wire net_U12043_Pad9;
    wire net_U12044_Pad10;
    wire net_U12044_Pad11;
    wire net_U12044_Pad9;
    wire net_U12045_Pad11;
    wire net_U12046_Pad6;
    wire net_U12046_Pad8;
    wire net_U12048_Pad6;
    wire net_U12049_Pad1;

    pullup R12001(__A12_1__GNZRO);
    pullup R12002(RELPLS);
    pullup R12003(INHPLS);
    pullup R12004(PALE);
    U74HC04 U12001(G01, __A12_1__G01A_n, G02, __A12_1__uG02_n, G03, __A12_1__uG03_n, GND, __A12_1__PA03_n, __A12_1__PA03, net_U12001_Pad10, G04, net_U12001_Pad12, G05, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12002(G01, G02, G01, __A12_1__uG02_n, __A12_1__uG03_n, net_U12002_Pad6, GND, net_U12002_Pad8, __A12_1__G01A_n, G02, __A12_1__uG03_n, net_U12002_Pad12, G03, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12003(__A12_1__G01A_n, __A12_1__uG02_n, G04, G05, G06, net_U12003_Pad6, GND, net_U12003_Pad8, G04, net_U12001_Pad12, net_U12003_Pad11, net_U12003_Pad12, G03, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12004(__A12_1__PA03, net_U12002_Pad12, net_U12002_Pad6, net_U12002_Pad8, net_U12003_Pad12,  , GND,  , net_U12003_Pad6, net_U12003_Pad8, net_U12004_Pad11, net_U12004_Pad12, __A12_1__PA06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12005(G06, net_U12003_Pad11, net_U12003_Pad6, net_U12005_Pad4, __A12_1__PA06, __A12_1__PA06_n, GND, net_U12005_Pad8, G07, net_U12005_Pad10, G08, net_U12005_Pad12, G09, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12006(net_U12001_Pad10, G05, net_U12001_Pad10, net_U12001_Pad12, G06, net_U12004_Pad12, GND, net_U12006_Pad8, G07, G08, G09, net_U12004_Pad11, net_U12003_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12007(G07, net_U12005_Pad10, net_U12005_Pad8, G08, net_U12005_Pad12, net_U12007_Pad6, GND, net_U12007_Pad8, net_U12005_Pad8, net_U12005_Pad10, G09, net_U12007_Pad12, net_U12005_Pad12, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12008(__A12_1__PA09, net_U12006_Pad8, net_U12007_Pad12, net_U12007_Pad6, net_U12007_Pad8,  , GND,  , net_U12008_Pad9, net_U12008_Pad10, net_U12008_Pad11, net_U12008_Pad12, __A12_1__PA12, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12009(net_U12006_Pad8, net_U12009_Pad2, __A12_1__PA09, __A12_1__PA09_n, G10, net_U12009_Pad6, GND, net_U12009_Pad8, G11, net_U12009_Pad10, G12, net_U12009_Pad12, net_U12008_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12010(G10, G11, G10, net_U12009_Pad8, net_U12009_Pad10, net_U12008_Pad10, GND, net_U12008_Pad11, net_U12009_Pad6, G11, net_U12009_Pad10, net_U12008_Pad9, G12, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12011(net_U12009_Pad6, net_U12009_Pad8, G13, G14, G16, net_U12011_Pad6, GND, net_U12011_Pad8, G13, net_U12011_Pad10, __A12_1__G16A_n, net_U12008_Pad12, G12, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12012(__A12_1__PA12, __A12_1__PA12_n, G13, net_U12012_Pad4, G14, net_U12011_Pad10, GND, __A12_1__G16A_n, G16, net_U12012_Pad10, net_U12011_Pad6, __A12_1__PA15_n, __A12_1__PA15, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12013(net_U12012_Pad4, G14, net_U12012_Pad4, net_U12011_Pad10, G16, net_U12013_Pad6, GND, net_U12013_Pad8, net_U12005_Pad4, net_U12009_Pad2, net_U12009_Pad12, net_U12013_Pad12, __A12_1__G16A_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U12014(__A12_1__PA15, net_U12011_Pad6, net_U12011_Pad8, net_U12013_Pad12, net_U12013_Pad6,  , GND,  , EXTPLS, RELPLS, INHPLS, net_U12014_Pad12, net_U12014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12015(net_U12015_Pad1, net_U12012_Pad10, G15, net_U12015_Pad4, TSUDO_n, __A12_1__T7PHS4_n, GND, __A12_1__uG02_n, G03, net_U12015_Pad10, G02, __A12_1__uG03_n, net_U12015_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U12016(net_U12013_Pad8, __A12_1__GNZRO, net_U12015_Pad1, __A12_1__GNZRO, net_U12016_Pad5, RELPLS, GND, RELPLS, net_U12015_Pad10, INHPLS, net_U12016_Pad11, INHPLS, net_U12015_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC04 U12017(__A12_1__GNZRO, net_U12017_Pad2, net_U12002_Pad6, net_U12017_Pad4, net_U12015_Pad4, net_U12017_Pad6, GND, GEQZRO_n, net_U12017_Pad9, net_U12017_Pad10, RAD, __A12_1__PB09_n, __A12_1__PB09, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12018(net_U12017_Pad4, net_U12017_Pad2, net_U12017_Pad2, net_U12017_Pad6, __A12_1__G01A_n, net_U12016_Pad5, GND, net_U12016_Pad11, net_U12017_Pad2, G01, net_U12017_Pad6, EXTPLS, net_U12017_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12019(net_U12017_Pad9, net_U12017_Pad2, G02, G01, G03,  , GND,  , net_U12019_Pad9, net_U12019_Pad10, net_U12019_Pad11, net_U12019_Pad12, __A12_1__PB09, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12020(net_U12014_Pad12, net_U12014_Pad13, T12A, RADRZ, net_U12014_Pad13, net_U12017_Pad10, GND, net_U12017_Pad10, net_U12014_Pad12, RADRG, __A12_1__PA12, __A12_1__PA15, net_U12020_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12021(__A12_1__PA03, __A12_1__PA06, __A12_1__PA03, __A12_1__PA06_n, __A12_1__PA09_n, net_U12019_Pad10, GND, net_U12019_Pad11, __A12_1__PA03_n, __A12_1__PA06, __A12_1__PA09_n, net_U12019_Pad9, __A12_1__PA09, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U12022(__A12_1__PA03_n, __A12_1__PA06_n, net_U12022_Pad3, MONPAR, SAP, net_U12022_Pad6, GND, net_U12022_Pad8, SCAD, net_U12022_Pad10, GOJAM, net_U12019_Pad12, __A12_1__PA09, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12023(net_U12023_Pad1, __A12_1__PA12_n, __A12_1__PA15_n, __A12_1__PB15, net_U12020_Pad13, net_U12023_Pad1, GND, __A12_1__PB09_n, __A12_1__PB15, net_U12023_Pad10, __A12_1__PB09, __A12_1__PB15_n, net_U12023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12024(__A12_1__PB15, __A12_1__PB15_n, __A12_1__PC15, PC15_n, __A12_1__PC15, MGP_n, GND, GEMP, PC15_n, MSP, net_U12022_Pad6,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12025(__A12_1__PC15, net_U12023_Pad10, net_U12023_Pad13, net_U12022_Pad3, CGG, net_U12022_Pad6, GND, __A12_1__PC15, net_U12022_Pad3, net_U12022_Pad10, PC15_n, net_U12022_Pad6, net_U12025_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12026(TPARG_n, n8XP5, T07_n, PHS4_n, FUTEXT, __A12_1__T7PHS4, GND, net_U12026_Pad8, XB0_n, T02_n, net_U12026_Pad11, net_U12026_Pad12, net_U12025_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U12027(net_U12022_Pad8, PALE, net_U12026_Pad12, PALE,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12028(G01ED, WEDOPG_n, WL08_n, net_U12028_Pad4, WL08_n, WSG_n, GND, net_U12028_Pad4, net_U12028_Pad13, net_U12028_Pad10, net_U12028_Pad10, CSG, net_U12028_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12029(net_U12028_Pad10, S08, net_U12028_Pad13, S08_n, net_U12029_Pad5, S09, GND, S09_n, net_U12029_Pad9, S10, net_U12029_Pad11, S10_n, net_U12029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12030(G02ED, WEDOPG_n, WL09_n, net_U12030_Pad4, WL09_n, WSG_n, GND, net_U12030_Pad4, net_U12029_Pad9, net_U12029_Pad5, net_U12029_Pad5, CSG, net_U12029_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12031(G03ED, WEDOPG_n, WL10_n, net_U12031_Pad4, WL10_n, WSG_n, GND, net_U12031_Pad4, net_U12029_Pad13, net_U12029_Pad11, net_U12029_Pad11, CSG, net_U12029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12032(G04ED, WEDOPG_n, WL11_n, net_U12032_Pad4, WL11_n, WSG_n, GND, net_U12032_Pad4, net_U12032_Pad13, net_U12032_Pad10, net_U12032_Pad10, CSG, net_U12032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12033(net_U12032_Pad10, S11, net_U12032_Pad13, S11_n, net_U12033_Pad5, S12, GND, S12_n, net_U12033_Pad9, S01, net_U12033_Pad11, S01_n, net_U12033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12034(G05ED, WEDOPG_n, WL12_n, net_U12034_Pad4, WL12_n, WSG_n, GND, EDOP_n, T12A, net_U12034_Pad10, net_U12033_Pad5, CSG, net_U12033_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U12035(G06ED, WEDOPG_n, WL13_n, G07ED, WEDOPG_n, WL14_n, GND, WL01_n, WSG_n, net_U12035_Pad10, net_U12035_Pad10, net_U12033_Pad13, net_U12033_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12036(net_U12033_Pad13, net_U12033_Pad11, CSG, net_U12036_Pad4, WL02_n, WSG_n, GND, net_U12036_Pad4, net_U12036_Pad13, net_U12036_Pad10, net_U12036_Pad10, CSG, net_U12036_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12037(net_U12036_Pad10, S02, net_U12036_Pad13, S02_n, net_U12037_Pad5, S03, GND, S03_n, net_U12037_Pad9, S04, net_U12037_Pad11, S04_n, net_U12037_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U12038(net_U12038_Pad1, WL03_n, WSG_n, net_U12037_Pad5, net_U12038_Pad1, net_U12037_Pad9, GND, net_U12037_Pad5, CSG, net_U12037_Pad9, WL04_n, WSG_n, net_U12038_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U12039(net_U12037_Pad11, net_U12038_Pad13, net_U12037_Pad13, net_U12037_Pad13, net_U12037_Pad11, CSG, GND, WL05_n, WSG_n, net_U12039_Pad10, net_U12039_Pad10, net_U12039_Pad12, net_U12039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12040(net_U12039_Pad12, net_U12039_Pad13, CSG, net_U12040_Pad4, WL06_n, WSG_n, GND, net_U12040_Pad4, net_U12040_Pad13, net_U12040_Pad10, net_U12040_Pad10, CSG, net_U12040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12041(net_U12039_Pad13, S05, net_U12039_Pad12, S05_n, net_U12040_Pad10, S06, GND, S06_n, net_U12040_Pad13, S07, net_U12041_Pad11, S07_n, net_U12041_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U12042(net_U12042_Pad1, WL07_n, WSG_n, net_U12041_Pad11, net_U12042_Pad1, net_U12041_Pad13, GND, net_U12041_Pad11, CSG, net_U12041_Pad13,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12043(__A12_1__T7PHS4, __A12_1__T7PHS4_n,  ,  , OCTAD2, net_U12026_Pad11, GND, GINH, net_U12043_Pad9, __A12_2__G01A, __A12_1__G01A_n,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12044( ,  ,  ,  ,  ,  , GND,  , net_U12044_Pad9, net_U12044_Pad10, net_U12044_Pad11, net_U12034_Pad10, net_U12043_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U12045( ,  ,  , CYR_n, net_U12026_Pad8, net_U12044_Pad9, GND, CYR_n, T12A, net_U12044_Pad9, net_U12045_Pad11, net_U12044_Pad10, SR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12046(net_U12026_Pad11, T02_n, net_U12026_Pad11, T02_n, XB2_n, net_U12046_Pad6, GND, net_U12046_Pad8, net_U12026_Pad11, T02_n, XB3_n, net_U12045_Pad11, XB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U12047(net_U12044_Pad10, SR_n, T12A, CYL_n, net_U12046_Pad6, net_U12044_Pad11, GND, CYL_n, T12A, net_U12044_Pad11, net_U12046_Pad8, net_U12034_Pad10, EDOP_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U12048(n8XP5, net_U12034_Pad4, SUMA16_n, SUMB16_n, __A12_1__G01A_n, net_U12048_Pad6, GND,  ,  ,  ,  , net_U12033_Pad5, net_U12033_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12049(net_U12049_Pad1, __A12_2__G01A, __A12_1__G16A_n, G16SW_n, net_U12049_Pad1, net_U12048_Pad6, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U12050(PALE, MPAL_n,  ,  ,  ,  ,  ,  ,  ,  ,  ,  ,  ,  , SIM_RST, SIM_CLK); //FPGA#OD:2
endmodule