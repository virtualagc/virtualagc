`timescale 1ns/1ps
`default_nettype none

module ch77_alarm_box(SIM_RST, SIM_CLK, p4VSW, GND, MDT01, MT01, MDT02, MT05, MDT03, MT12, MDT04, MWL01, MDT05, MWL02, MDT06, MWL03, MDT07, MWL04, MDT08, MWL05, MDT09, MWL06, MDT10, MRCH, MDT11, MWCH, MDT12, MWSG, MDT13, MPAL_n, MDT14, MTCAL_n, MDT15, MRPTAL_n, MDT16, MWATCH_n, MNHSBF, MVFAIL_n, MNHNC, MCTRAL_n, MNHRPT, MSCAFL_n, MTCSAI, MSCDBL_n, MSTRT, MAMU, MSTP, MSBSTP, MRDCH, MLDCH, MONPAR, MONWBK, MLOAD, MREAD, NHALGA, DOSCAL, DBLTST);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    output wire DBLTST;
    output wire DOSCAL;
    output wire MAMU;
    input wire MCTRAL_n;
    output wire MDT01;
    output wire MDT02;
    output wire MDT03;
    output wire MDT04;
    output wire MDT05;
    output wire MDT06;
    output wire MDT07;
    output wire MDT08;
    output wire MDT09;
    output wire MDT10;
    output wire MDT11;
    output wire MDT12;
    output wire MDT13;
    output wire MDT14;
    output wire MDT15;
    output wire MDT16;
    output wire MLDCH;
    output wire MLOAD;
    output wire MNHNC;
    output wire MNHRPT;
    output wire MNHSBF;
    output wire MONPAR;
    output wire MONWBK;
    input wire MPAL_n;
    input wire MRCH;
    output wire MRDCH;
    output wire MREAD;
    input wire MRPTAL_n;
    output wire MSBSTP;
    input wire MSCAFL_n;
    input wire MSCDBL_n;
    output wire MSTP;
    output wire MSTRT;
    input wire MT01;
    input wire MT05;
    input wire MT12;
    input wire MTCAL_n;
    output wire MTCSAI;
    input wire MVFAIL_n;
    input wire MWATCH_n;
    input wire MWCH;
    input wire MWL01;
    input wire MWL02;
    input wire MWL03;
    input wire MWL04;
    input wire MWL05;
    input wire MWL06;
    input wire MWSG;
    output wire NHALGA;
    wire __RestartMonitor__CCH77;
    wire __RestartMonitor__RCH77_n;
    wire net_R77009_Pad2; //FPGA#wand
    wire net_U77001_Pad10;
    wire net_U77001_Pad12;
    wire net_U77001_Pad2;
    wire net_U77001_Pad4;
    wire net_U77001_Pad6;
    wire net_U77001_Pad8;
    wire net_U77002_Pad11;
    wire net_U77002_Pad12;
    wire net_U77002_Pad2;
    wire net_U77002_Pad4;
    wire net_U77002_Pad6;
    wire net_U77002_Pad8;
    wire net_U77003_Pad1;
    wire net_U77003_Pad13;
    wire net_U77005_Pad1;
    wire net_U77005_Pad12;
    wire net_U77006_Pad1;
    wire net_U77006_Pad10;
    wire net_U77006_Pad13;
    wire net_U77006_Pad3;
    wire net_U77006_Pad8;
    wire net_U77007_Pad10;
    wire net_U77007_Pad11;
    wire net_U77007_Pad12;
    wire net_U77007_Pad13;
    wire net_U77007_Pad3;
    wire net_U77007_Pad4;
    wire net_U77007_Pad5;
    wire net_U77008_Pad10;
    wire net_U77008_Pad12;
    wire net_U77008_Pad8;
    wire net_U77009_Pad10;
    wire net_U77009_Pad12;
    wire net_U77009_Pad13;
    wire net_U77009_Pad4;
    wire net_U77010_Pad10;
    wire net_U77010_Pad11;
    wire net_U77010_Pad12;
    wire net_U77010_Pad13;
    wire net_U77010_Pad4;
    wire net_U77011_Pad10;
    wire net_U77011_Pad4;
    wire net_U77011_Pad5;

    pullup R77001(MWL01);
    pullup R77002(MWL02);
    pullup R77003(MWL03);
    pullup R77004(MWL04);
    pullup R77005(MWL05);
    pullup R77006(MWL06);
    pullup R77007(MT01);
    pullup R77008(MWSG);
    pullup R77009(net_R77009_Pad2);
    pullup R77010(MT12);
    pullup R77011(MWCH);
    pullup R77012(MRCH);
    pullup R77013(MT05);
    pullup R77014(MTCAL_n);
    pullup R77015(MRPTAL_n);
    pullup R77016(MWATCH_n);
    pullup R77017(MVFAIL_n);
    pullup R77018(MCTRAL_n);
    pullup R77019(MSCAFL_n);
    pullup R77020(MSCDBL_n);
    pulldown R77021(MDT10);
    pulldown R77022(MDT11);
    pulldown R77023(MDT12);
    pulldown R77024(MDT13);
    pulldown R77025(MDT14);
    pulldown R77026(MDT15);
    pulldown R77027(MDT16);
    pulldown R77028(MNHSBF);
    pulldown R77029(MNHNC);
    pulldown R77030(MNHRPT);
    pulldown R77031(MTCSAI);
    pulldown R77032(MSTRT);
    pulldown R77033(MSTP);
    pulldown R77034(MSBSTP);
    pulldown R77035(MRDCH);
    pulldown R77036(MLDCH);
    pulldown R77037(MONPAR);
    pulldown R77038(MONWBK);
    pulldown R77039(MLOAD);
    pulldown R77040(MREAD);
    pulldown R77041(NHALGA);
    pulldown R77042(DOSCAL);
    pulldown R77043(DBLTST);
    pulldown R77044(MAMU);
    pullup R77045(MPAL_n);
    U74HC04 U77001(MWL01, net_U77001_Pad2, MWL02, net_U77001_Pad4, MWL03, net_U77001_Pad6, GND, net_U77001_Pad8, MWL04, net_U77001_Pad10, MWL05, net_U77001_Pad12, MWL06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0) U77002(MT01, net_U77002_Pad2, MWSG, net_U77002_Pad4, MWCH, net_U77002_Pad6, GND, net_U77002_Pad8, MRCH, __RestartMonitor__RCH77_n, net_U77002_Pad11, net_U77002_Pad12, MPAL_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U77003(net_U77003_Pad1, net_U77001_Pad2, net_U77001_Pad4, net_U77001_Pad6, net_U77001_Pad8,  , GND,  , net_U77001_Pad10, net_U77001_Pad12, net_U77002_Pad2, net_U77002_Pad4, net_U77003_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U77004(net_U77003_Pad1, net_R77009_Pad2, net_U77003_Pad13, net_R77009_Pad2,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U77005(net_U77005_Pad1, MT12, net_U77005_Pad12, net_U77005_Pad12, net_U77005_Pad1, net_R77009_Pad2, GND, net_U77002_Pad8, net_U77005_Pad12, net_U77002_Pad11, net_U77002_Pad6, net_U77005_Pad12, __RestartMonitor__CCH77, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U77006(net_U77006_Pad1, net_U77002_Pad12, net_U77006_Pad3, net_U77006_Pad3, net_U77006_Pad1, __RestartMonitor__CCH77, GND, net_U77006_Pad8, net_U77006_Pad13, net_U77006_Pad10, net_U77006_Pad10, __RestartMonitor__CCH77, net_U77006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U77007(net_U77006_Pad8, MPAL_n, net_U77007_Pad3, net_U77007_Pad4, net_U77007_Pad5, net_U77007_Pad10, GND, net_U77007_Pad4, __RestartMonitor__CCH77, net_U77007_Pad10, net_U77007_Pad11, net_U77007_Pad12, net_U77007_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U77008(MT05, net_U77007_Pad3, MTCAL_n, net_U77007_Pad5, MRPTAL_n, net_U77007_Pad11, GND, net_U77008_Pad8, MWATCH_n, net_U77008_Pad10, MVFAIL_n, net_U77008_Pad12, MCTRAL_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U77009(net_U77007_Pad12, net_U77007_Pad13, __RestartMonitor__CCH77, net_U77009_Pad4, net_U77008_Pad8, net_U77009_Pad10, GND, net_U77009_Pad4, __RestartMonitor__CCH77, net_U77009_Pad10, net_U77008_Pad10, net_U77009_Pad12, net_U77009_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U77010(net_U77009_Pad12, net_U77009_Pad13, __RestartMonitor__CCH77, net_U77010_Pad4, net_U77008_Pad12, net_U77010_Pad10, GND, net_U77010_Pad4, __RestartMonitor__CCH77, net_U77010_Pad10, net_U77010_Pad11, net_U77010_Pad12, net_U77010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U77011(net_U77010_Pad12, net_U77010_Pad13, __RestartMonitor__CCH77, net_U77011_Pad4, net_U77011_Pad5, net_U77011_Pad10, GND, net_U77011_Pad4, __RestartMonitor__CCH77, net_U77011_Pad10,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U77012(MSCAFL_n, net_U77010_Pad11, MSCDBL_n, net_U77011_Pad5,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U77013(__RestartMonitor__RCH77_n, net_U77006_Pad1, __RestartMonitor__RCH77_n, net_U77006_Pad10, GND, MDT02, GND, MDT03, __RestartMonitor__RCH77_n, net_U77007_Pad4, GND, MDT01, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U77014(__RestartMonitor__RCH77_n, net_U77007_Pad13, __RestartMonitor__RCH77_n, net_U77009_Pad4, GND, MDT05, GND, MDT06, __RestartMonitor__RCH77_n, net_U77009_Pad13, GND, MDT04, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U77015(__RestartMonitor__RCH77_n, net_U77010_Pad4, __RestartMonitor__RCH77_n, net_U77010_Pad13, GND, MDT08, GND, MDT09, __RestartMonitor__RCH77_n, net_U77011_Pad4, GND, MDT07, GND, p4VSW, SIM_RST, SIM_CLK);
endmodule