// Verilog testbench created by dumbTestbench.py
`timescale 100ns / 1ns

module agc;

reg rst = 1;
reg STRT2 = 1;
initial
  begin
    $dumpfile("agc.lxt2");
    $dumpvars(0, agc);
    # 1 rst = 0;
    # 50 STRT2 = 0;
    # 1000 $finish;
  end

reg CLOCK = 0;
always #2.44140625 CLOCK = !CLOCK;

reg ALTEST = 0, CAURST = 0, CCH13 = 0, CCH33 = 0, CGA18 = 0, CH1111 = 0,
  CH1112 = 0, CH1114 = 0, CH1116 = 0, CH1211 = 0, CH1212 = 0, CH1216 = 0,
  CH3311 = 0, CH3313 = 0, CH3314 = 0, CH3316 = 0, CHAT11 = 0, CHAT12 = 0,
  CHAT13 = 0, CHAT14 = 0, CHBT11 = 0, CHBT12 = 0, CHBT13 = 0, CHBT14 = 0,
  CHOR11_ = 0, CHOR12_ = 0, CHOR13_ = 0, CHOR16_ = 0, CHWL01_ = 0, CHWL02_ = 0,
  CHWL03_ = 0, CHWL04_ = 0, CHWL11_ = 0, DKEND = 0, F09A_ = 0, F09B = 0,
  F09B_ = 0, F09D = 0, F10A = 0, F10A_ = 0, F17A = 0, F17B = 0, F5ASB2_ = 0,
  F5BSB2_ = 0, GOJAM = 0, GTRST_ = 0, GTSET_ = 0, LRIN0 = 0, LRIN1 = 0,
  MAINRS = 0, MARK = 0, MKEY1 = 0, MKEY2 = 0, MKEY3 = 0, MKEY4 = 0, MKEY5 = 0,
  MRKREJ = 0, MRKRST = 0, NAVRST = 0, NKEY1 = 0, NKEY2 = 0, NKEY3 = 0,
  NKEY4 = 0, NKEY5 = 0, RCH13_ = 0, RCH33_ = 0, RCHG_ = 0, RRIN0 = 0, RRIN1 = 0,
  SB0_ = 0, SB2_ = 0, SBYBUT = 0, STOP = 0, T05 = 0, T11 = 0, TEMPIN = 0,
  W1110 = 0, WCH13_ = 0, XB5_ = 0, XB6_ = 0, XT1_ = 0;

wire CH11, CH12, CH13, CH1301, CH1302, CH1303, CH1304, CH1311, CH14, CH1501,
  CH1502, CH1503, CH1504, CH1505, CH16, CH1601, CH1602, CH1603, CH1604,
  CH1605, CH1606, CH1607, CH3312, CHOR14_, CNTOF9, DLKRPT, END, ERRST,
  F10AS0, F17A_, F17B_, HERB, KYRPT1, KYRPT2, LRRANG, LRSYNC, LRXVEL, LRYVEL,
  LRZVEL, MKRPT, RADRPT, RCH15_, RCH16_, RNRADM, RNRADP, RRRANG, RRRARA,
  RRSYNC, SBY, SBYLIT, STNDBY, STNDBY_, TEMPIN_, TPORA_, TPOR_;

A18 iA18 (
  rst, ALTEST, CAURST, CCH13, CCH33, CGA18, CH1111, CH1112, CH1114, CH1116,
  CH1211, CH1212, CH1216, CH3311, CH3313, CH3314, CH3316, CHAT11, CHAT12,
  CHAT13, CHAT14, CHBT11, CHBT12, CHBT13, CHBT14, CHOR11_, CHOR12_, CHOR13_,
  CHOR16_, CHWL01_, CHWL02_, CHWL03_, CHWL04_, CHWL11_, DKEND, F09A_, F09B,
  F09B_, F09D, F10A, F10A_, F17A, F17B, F5ASB2_, F5BSB2_, GOJAM, GTRST_,
  GTSET_, LRIN0, LRIN1, MAINRS, MARK, MKEY1, MKEY2, MKEY3, MKEY4, MKEY5,
  MRKREJ, MRKRST, NAVRST, NKEY1, NKEY2, NKEY3, NKEY4, NKEY5, RCH13_, RCH33_,
  RCHG_, RRIN0, RRIN1, SB0_, SB2_, SBYBUT, STOP, T05, T11, TEMPIN, W1110,
  WCH13_, XB5_, XB6_, XT1_, CHOR14_, F17A_, F17B_, HERB, TPORA_, TPOR_, CH11,
  CH12, CH13, CH1301, CH1302, CH1303, CH1304, CH1311, CH14, CH1501, CH1502,
  CH1503, CH1504, CH1505, CH16, CH1601, CH1602, CH1603, CH1604, CH1605, CH1606,
  CH1607, CH3312, CNTOF9, DLKRPT, END, ERRST, F10AS0, KYRPT1, KYRPT2, LRRANG,
  LRSYNC, LRXVEL, LRYVEL, LRZVEL, MKRPT, RADRPT, RCH15_, RCH16_, RNRADM,
  RNRADP, RRRANG, RRRARA, RRSYNC, SBY, SBYLIT, STNDBY, STNDBY_, TEMPIN_
);

initial $timeformat(-9, 0, " ns", 10);
initial $monitor("%t: %d", $time, CLOCK);

endmodule
