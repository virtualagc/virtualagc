`timescale 1ns/1ps
`default_nettype none

module inout_ii(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, F04B, FS05_n, F05A_n, F05B_n, TPOR_n, CCHG_n, WCHG_n, IN3301, ULLTHR, RRPONA, SMSEPR, RRRLSC, SPSRDY, ZEROP, S4BSAB, OPMSW2, LFTOFF, OPMSW3, GUIREL, STRPRS, OPCDFL, LVDAGD, IN3008, LRRLSC, IMUOPR, CH3310, CTLSAT, LEMATT, IMUCAG, IN3212, CDUFAL, HOLFUN, IN3213, IMUFAL, FREFUN, IN3214, ISSTOR, GCAPCL, IN3216, TEMPIN, TRST9, TRST10, PCHGOF, ROLGOF, MANpP, MANmP, MANpY, MANmY, MANpR, MANmR, TRANpX, TRANmX, TRANpY, TRANmY, TRANpZ, TRANmZ, MNIMpP, MNIMmP, MNIMpY, MNIMmY, MNIMpR, MNIMmR, PIPAFL, AGCWAR, OSCALM, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CHWL16_n, CH1213, CH1214, CH1301, CH1302, CH1303, CH1304, CH1305, CH1306, CH1307, CH1308, CH1309, CH1310, CH1311, CH1316, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406, CH1407, CH1408, CH1409, CH1410, CH1411, CH1412, CH1413, CH1414, CH1416, CH3312, XB0_n, XB1_n, XB2_n, XB3_n, XT1_n, XT3_n, WCH13_n, CCH11, RCH11_n, RCH33_n, WCH11_n, HNDRPT, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207, CH3208, CH3209, CH3210, CH3313, CH3314, CH3316, CHOR01_n, CHOR02_n, CHOR03_n, CHOR04_n, CHOR05_n, CHOR06_n, CHOR07_n, CHOR08_n, CHOR09_n, CHOR10_n, CHOR11_n, CHOR12_n, CHOR13_n, CHOR14_n, CHOR16_n, RLYB01, RLYB02, RLYB03, RLYB04, RLYB05, RLYB06, RLYB07, RLYB08, RLYB09, RLYB10, RLYB11, RYWD12, RYWD13, RYWD14, RYWD16);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire AGCWAR;
    output wire CCH11;
    input wire CCHG_n;
    input wire CDUFAL;
    input wire CH1213;
    input wire CH1214;
    input wire CH1301;
    input wire CH1302;
    input wire CH1303;
    input wire CH1304;
    input wire CH1305;
    input wire CH1306;
    input wire CH1307;
    input wire CH1308;
    input wire CH1309;
    input wire CH1310;
    input wire CH1311;
    input wire CH1316;
    input wire CH1401;
    input wire CH1402;
    input wire CH1403;
    input wire CH1404;
    input wire CH1405;
    input wire CH1406;
    input wire CH1407;
    input wire CH1408;
    input wire CH1409;
    input wire CH1410;
    input wire CH1411;
    input wire CH1412;
    input wire CH1413;
    input wire CH1414;
    input wire CH1416;
    output wire CH3201;
    output wire CH3202;
    output wire CH3203;
    output wire CH3204;
    output wire CH3205;
    output wire CH3206;
    output wire CH3207;
    output wire CH3208;
    output wire CH3209;
    output wire CH3210;
    input wire CH3310;
    input wire CH3312;
    output wire CH3313;
    output wire CH3314;
    output wire CH3316;
    output wire CHOR01_n; //FPGA#wand
    output wire CHOR02_n; //FPGA#wand
    output wire CHOR03_n; //FPGA#wand
    output wire CHOR04_n; //FPGA#wand
    output wire CHOR05_n; //FPGA#wand
    output wire CHOR06_n; //FPGA#wand
    output wire CHOR07_n; //FPGA#wand
    output wire CHOR08_n; //FPGA#wand
    output wire CHOR09_n; //FPGA#wand
    output wire CHOR10_n; //FPGA#wand
    output wire CHOR11_n; //FPGA#wand
    output wire CHOR12_n; //FPGA#wand
    output wire CHOR13_n; //FPGA#wand
    output wire CHOR14_n; //FPGA#wand
    output wire CHOR16_n; //FPGA#wand
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire CHWL16_n;
    input wire CTLSAT;
    input wire F04B;
    input wire F05A_n;
    input wire F05B_n;
    input wire FREFUN;
    input wire FS05_n;
    input wire GCAPCL;
    input wire GOJAM;
    input wire GUIREL;
    output wire HNDRPT;
    input wire HOLFUN;
    input wire IMUCAG;
    input wire IMUFAL;
    input wire IMUOPR;
    input wire IN3008;
    input wire IN3212;
    input wire IN3213;
    input wire IN3214;
    input wire IN3216;
    input wire IN3301;
    input wire ISSTOR;
    input wire LEMATT;
    input wire LFTOFF;
    input wire LRRLSC;
    input wire LVDAGD;
    input wire MANmP;
    input wire MANmR;
    input wire MANmY;
    input wire MANpP;
    input wire MANpR;
    input wire MANpY;
    input wire MNIMmP;
    input wire MNIMmR;
    input wire MNIMmY;
    input wire MNIMpP;
    input wire MNIMpR;
    input wire MNIMpY;
    input wire OPCDFL;
    input wire OPMSW2;
    input wire OPMSW3;
    input wire OSCALM;
    input wire PCHGOF;
    input wire PIPAFL;
    output wire RCH11_n;
    output wire RCH33_n;
    output wire RLYB01;
    output wire RLYB02;
    output wire RLYB03;
    output wire RLYB04;
    output wire RLYB05;
    output wire RLYB06;
    output wire RLYB07;
    output wire RLYB08;
    output wire RLYB09;
    output wire RLYB10;
    output wire RLYB11;
    input wire ROLGOF;
    input wire RRPONA;
    input wire RRRLSC;
    output wire RYWD12;
    output wire RYWD13;
    output wire RYWD14;
    output wire RYWD16;
    input wire S4BSAB;
    input wire SMSEPR;
    input wire SPSRDY;
    input wire STRPRS;
    input wire TEMPIN;
    input wire TPOR_n;
    input wire TRANmX;
    input wire TRANmY;
    input wire TRANmZ;
    input wire TRANpX;
    input wire TRANpY;
    input wire TRANpZ;
    input wire TRST10;
    input wire TRST9;
    input wire ULLTHR;
    output wire WCH11_n;
    input wire WCH13_n;
    input wire WCHG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    input wire XT1_n;
    input wire XT3_n;
    input wire ZEROP;
    wire __A17_1__F04B_n;
    wire __A17_1__FO5D;
    wire __A17_1__RCH30_n;
    wire __A17_1__RCH31_n;
    wire __A17_1__RCH32_n;
    wire __A17_1__TRP31A;
    wire __A17_1__TRP31B;
    wire __A17_1__TRP32;
    wire __A17_2__CCH10;
    wire __A17_2__RCH10_n;
    wire __A17_2__WCH10_n;
    wire net_R17016_Pad2; //FPGA#wand
    wire net_R17017_Pad2; //FPGA#wand
    wire net_R17018_Pad2; //FPGA#wand
    wire net_U17001_Pad1;
    wire net_U17001_Pad10;
    wire net_U17001_Pad13;
    wire net_U17001_Pad4;
    wire net_U17002_Pad13;
    wire net_U17002_Pad5;
    wire net_U17002_Pad9;
    wire net_U17003_Pad1;
    wire net_U17003_Pad11;
    wire net_U17003_Pad13;
    wire net_U17003_Pad3;
    wire net_U17003_Pad5;
    wire net_U17003_Pad9;
    wire net_U17004_Pad1;
    wire net_U17004_Pad10;
    wire net_U17004_Pad13;
    wire net_U17005_Pad1;
    wire net_U17005_Pad10;
    wire net_U17005_Pad13;
    wire net_U17005_Pad4;
    wire net_U17007_Pad1;
    wire net_U17007_Pad10;
    wire net_U17007_Pad13;
    wire net_U17007_Pad4;
    wire net_U17008_Pad10;
    wire net_U17008_Pad11;
    wire net_U17008_Pad3;
    wire net_U17008_Pad5;
    wire net_U17008_Pad9;
    wire net_U17010_Pad10;
    wire net_U17010_Pad13;
    wire net_U17010_Pad4;
    wire net_U17011_Pad10;
    wire net_U17011_Pad11;
    wire net_U17011_Pad12;
    wire net_U17011_Pad3;
    wire net_U17011_Pad4;
    wire net_U17011_Pad5;
    wire net_U17011_Pad6;
    wire net_U17011_Pad8;
    wire net_U17011_Pad9;
    wire net_U17012_Pad11;
    wire net_U17012_Pad13;
    wire net_U17012_Pad9;
    wire net_U17014_Pad10;
    wire net_U17014_Pad13;
    wire net_U17015_Pad10;
    wire net_U17015_Pad11;
    wire net_U17015_Pad3;
    wire net_U17015_Pad4;
    wire net_U17015_Pad5;
    wire net_U17015_Pad9;
    wire net_U17017_Pad10;
    wire net_U17017_Pad13;
    wire net_U17018_Pad10;
    wire net_U17018_Pad11;
    wire net_U17018_Pad12;
    wire net_U17018_Pad13;
    wire net_U17018_Pad3;
    wire net_U17018_Pad4;
    wire net_U17018_Pad5;
    wire net_U17018_Pad6;
    wire net_U17018_Pad8;
    wire net_U17018_Pad9;
    wire net_U17019_Pad11;
    wire net_U17019_Pad13;
    wire net_U17019_Pad9;
    wire net_U17022_Pad8;
    wire net_U17022_Pad9;
    wire net_U17023_Pad1;
    wire net_U17023_Pad10;
    wire net_U17023_Pad6;
    wire net_U17023_Pad9;
    wire net_U17025_Pad10;
    wire net_U17025_Pad11;
    wire net_U17025_Pad5;
    wire net_U17025_Pad6;
    wire net_U17026_Pad12;
    wire net_U17026_Pad3;
    wire net_U17027_Pad11;
    wire net_U17027_Pad13;
    wire net_U17027_Pad3;
    wire net_U17027_Pad5;
    wire net_U17027_Pad9;
    wire net_U17028_Pad12;
    wire net_U17031_Pad11;
    wire net_U17031_Pad12;
    wire net_U17031_Pad13;
    wire net_U17033_Pad12;
    wire net_U17033_Pad3;
    wire net_U17034_Pad11;
    wire net_U17034_Pad4;
    wire net_U17034_Pad9;
    wire net_U17035_Pad10;
    wire net_U17036_Pad13;
    wire net_U17037_Pad13;
    wire net_U17037_Pad3;
    wire net_U17038_Pad1;
    wire net_U17038_Pad10;
    wire net_U17038_Pad13;
    wire net_U17038_Pad3;
    wire net_U17039_Pad11;
    wire net_U17039_Pad13;
    wire net_U17039_Pad3;
    wire net_U17039_Pad5;
    wire net_U17039_Pad9;
    wire net_U17040_Pad10;
    wire net_U17040_Pad12;
    wire net_U17040_Pad4;
    wire net_U17040_Pad6;
    wire net_U17040_Pad8;
    wire net_U17041_Pad11;
    wire net_U17041_Pad13;
    wire net_U17041_Pad9;
    wire net_U17042_Pad13;
    wire net_U17042_Pad3;
    wire net_U17043_Pad13;
    wire net_U17043_Pad3;
    wire net_U17044_Pad10;
    wire net_U17044_Pad13;
    wire net_U17044_Pad3;
    wire net_U17045_Pad4;
    wire net_U17046_Pad13;
    wire net_U17046_Pad3;
    wire net_U17047_Pad10;
    wire net_U17047_Pad13;
    wire net_U17047_Pad3;
    wire net_U17048_Pad10;
    wire net_U17048_Pad4;
    wire net_U17048_Pad8;
    wire net_U17049_Pad1;
    wire net_U17049_Pad13;
    wire net_U17049_Pad3;
    wire net_U17050_Pad11;
    wire net_U17050_Pad13;
    wire net_U17050_Pad3;
    wire net_U17050_Pad5;
    wire net_U17050_Pad9;
    wire net_U17051_Pad13;
    wire net_U17051_Pad3;
    wire net_U17052_Pad11;
    wire net_U17052_Pad13;
    wire net_U17052_Pad3;
    wire net_U17052_Pad5;
    wire net_U17052_Pad9;
    wire net_U17053_Pad10;
    wire net_U17053_Pad13;
    wire net_U17053_Pad3;
    wire net_U17054_Pad10;
    wire net_U17054_Pad4;
    wire net_U17055_Pad13;
    wire net_U17055_Pad3;
    wire net_U17056_Pad13;
    wire net_U17056_Pad3;
    wire net_U17057_Pad10;
    wire net_U17057_Pad13;
    wire net_U17057_Pad3;
    wire net_U17058_Pad1;
    wire net_U17058_Pad10;
    wire net_U17058_Pad13;
    wire net_U17058_Pad3;
    wire net_U17059_Pad13;
    wire net_U17059_Pad3;
    wire net_U17059_Pad5;
    wire net_U17059_Pad9;
    wire net_U17060_Pad10;
    wire net_U17060_Pad11;
    wire net_U17060_Pad3;
    wire net_U17061_Pad1;
    wire net_U17063_Pad8;
    wire net_U17064_Pad1;
    wire net_U17064_Pad10;

    pullup R17001(CHOR01_n);
    pullup R17002(CHOR02_n);
    pullup R17003(CHOR03_n);
    pullup R17004(CHOR04_n);
    pullup R17005(CHOR05_n);
    pullup R17006(CHOR06_n);
    pullup R17007(CHOR07_n);
    pullup R17008(CHOR08_n);
    pullup R17009(CHOR09_n);
    pullup R17010(CHOR10_n);
    pullup R17011(CHOR11_n);
    pullup R17012(CHOR12_n);
    pullup R17013(CHOR13_n);
    pullup R17014(CHOR14_n);
    pullup R17015(CHOR16_n);
    pullup R17016(net_R17016_Pad2);
    pullup R17017(net_R17017_Pad2);
    pullup R17018(net_R17018_Pad2);
    U74HC02 U17001(net_U17001_Pad1, IN3301, RCH33_n, net_U17001_Pad4, XB3_n, XT3_n, GND, ULLTHR, __A17_1__RCH30_n, net_U17001_Pad10, XB0_n, XT3_n, net_U17001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17002(net_U17001_Pad4, RCH33_n, net_U17001_Pad13, __A17_1__RCH30_n, net_U17002_Pad5, __A17_1__RCH31_n, GND, __A17_1__RCH32_n, net_U17002_Pad9, __A17_1__F04B_n, F04B, RLYB01, net_U17002_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17003(net_U17003_Pad1, CHOR01_n, net_U17003_Pad3, CHOR02_n, net_U17003_Pad5, CHOR03_n, GND, CHOR04_n, net_U17003_Pad9, CHOR05_n, net_U17003_Pad11, CHOR06_n, net_U17003_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U17004(net_U17004_Pad1, MANpP, __A17_1__RCH31_n, net_U17002_Pad5, XB1_n, XT3_n, GND, SMSEPR, __A17_1__RCH30_n, net_U17004_Pad10, RRPONA, RCH33_n, net_U17004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17005(net_U17005_Pad1, MANmP, __A17_1__RCH31_n, net_U17005_Pad4, RRRLSC, RCH33_n, GND, MANpY, __A17_1__RCH31_n, net_U17005_Pad10, SPSRDY, __A17_1__RCH30_n, net_U17005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17006(net_U17001_Pad1, net_U17001_Pad10, net_U17004_Pad13, net_U17004_Pad10, net_U17005_Pad1, net_U17003_Pad3, GND, net_U17003_Pad5, net_U17005_Pad4, net_U17005_Pad13, net_U17005_Pad10, net_U17003_Pad1, net_U17004_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17007(net_U17007_Pad1, S4BSAB, __A17_1__RCH30_n, net_U17007_Pad4, ZEROP, RCH33_n, GND, MANmY, __A17_1__RCH31_n, net_U17007_Pad10, LFTOFF, __A17_1__RCH30_n, net_U17007_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17008(net_U17007_Pad4, net_U17007_Pad1, net_U17008_Pad3, net_U17007_Pad13, net_U17008_Pad5, net_U17003_Pad11, GND, net_U17003_Pad13, net_U17008_Pad9, net_U17008_Pad10, net_U17008_Pad11, net_U17003_Pad9, net_U17007_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17009(net_U17008_Pad3, OPMSW2, RCH33_n, net_U17008_Pad5, MANpR, __A17_1__RCH31_n, GND, GUIREL, __A17_1__RCH30_n, net_U17008_Pad10, OPMSW3, RCH33_n, net_U17008_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17010(net_U17008_Pad11, MANmR, __A17_1__RCH31_n, net_U17010_Pad4, OPCDFL, __A17_1__RCH30_n, GND, STRPRS, RCH33_n, net_U17010_Pad10, TRANpX, __A17_1__RCH31_n, net_U17010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17011(net_U17010_Pad10, net_U17010_Pad4, net_U17011_Pad3, net_U17011_Pad4, net_U17011_Pad5, net_U17011_Pad6, GND, net_U17011_Pad8, net_U17011_Pad9, net_U17011_Pad10, net_U17011_Pad11, net_U17011_Pad12, net_U17010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17012(net_U17011_Pad12, CHOR07_n, net_U17011_Pad6, CHOR08_n, net_U17011_Pad8, CHOR09_n, GND, CHOR10_n, net_U17012_Pad9, CHOR11_n, net_U17012_Pad11, CHOR12_n, net_U17012_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U17013(net_U17011_Pad4, IN3008, __A17_1__RCH30_n, net_U17011_Pad3, LVDAGD, RCH33_n, GND, TRANmX, __A17_1__RCH31_n, net_U17011_Pad5, IMUOPR, __A17_1__RCH30_n, net_U17011_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17014(net_U17011_Pad9, LRRLSC, RCH33_n, net_U17011_Pad11, TRANpY, __A17_1__RCH31_n, GND, CTLSAT, __A17_1__RCH30_n, net_U17014_Pad10, TRANmY, __A17_1__RCH31_n, net_U17014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17015(CH3310, net_U17014_Pad10, net_U17015_Pad3, net_U17015_Pad4, net_U17015_Pad5, net_U17012_Pad11, GND, net_U17012_Pad13, net_U17015_Pad9, net_U17015_Pad10, net_U17015_Pad11, net_U17012_Pad9, net_U17014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17016(net_U17015_Pad4, IMUCAG, __A17_1__RCH30_n, net_U17015_Pad3, LEMATT, __A17_1__RCH32_n, GND, TRANpZ, __A17_1__RCH31_n, net_U17015_Pad5, CDUFAL, __A17_1__RCH30_n, net_U17015_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17017(net_U17015_Pad9, IN3212, __A17_1__RCH32_n, net_U17015_Pad11, TRANmZ, __A17_1__RCH31_n, GND, IMUFAL, __A17_1__RCH30_n, net_U17017_Pad10, IN3213, __A17_1__RCH32_n, net_U17017_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17018(net_U17017_Pad13, net_U17017_Pad10, net_U17018_Pad3, net_U17018_Pad4, net_U17018_Pad5, net_U17018_Pad6, GND, net_U17018_Pad8, net_U17018_Pad9, net_U17018_Pad10, net_U17018_Pad11, net_U17018_Pad12, net_U17018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17019(net_U17018_Pad12, CHOR13_n, net_U17018_Pad6, CHOR14_n, net_U17018_Pad8, CHOR16_n, GND, net_R17016_Pad2, net_U17019_Pad9, net_R17016_Pad2, net_U17019_Pad11, net_R17017_Pad2, net_U17019_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U17020(net_U17018_Pad13, HOLFUN, __A17_1__RCH31_n, net_U17018_Pad4, ISSTOR, __A17_1__RCH30_n, GND, IN3214, __A17_1__RCH32_n, net_U17018_Pad3, FREFUN, __A17_1__RCH31_n, net_U17018_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17021(net_U17018_Pad10, TEMPIN, __A17_1__RCH30_n, net_U17018_Pad9, IN3216, __A17_1__RCH32_n, GND, GCAPCL, __A17_1__RCH31_n, net_U17018_Pad11, XB2_n, XT3_n, net_U17002_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17022(MANpP, MANmP, MANmY, MANpR, MANmR, net_U17019_Pad11, GND, net_U17022_Pad8, net_U17022_Pad9, net_R17016_Pad2, F05A_n, net_U17019_Pad9, MANpY, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U17023(net_U17023_Pad1, CHWL12_n, WCH13_n, net_U17022_Pad9, net_U17023_Pad1, net_U17023_Pad6, GND, net_U17022_Pad8, net_U17023_Pad9, net_U17023_Pad10, __A17_1__F04B_n, FS05_n, __A17_1__FO5D, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17024(net_U17022_Pad9, GOJAM, net_U17023_Pad10, net_R17016_Pad2, __A17_1__FO5D, net_U17023_Pad9, GND, net_U17019_Pad13, TRANpX, TRANmX, TRANpY, net_U17023_Pad6, __A17_1__TRP31A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U17025(__A17_1__TRP31A, net_U17023_Pad10, F05B_n, net_U17025_Pad11, net_U17025_Pad5, net_U17025_Pad6, GND, CHWL13_n, WCH13_n, net_U17025_Pad10, net_U17025_Pad11, F05B_n, __A17_1__TRP31B, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17026(TRANmY, TRANpZ, net_U17026_Pad3, net_R17017_Pad2, F05A_n, net_U17025_Pad5, GND, net_U17025_Pad6, net_U17025_Pad11, net_R17017_Pad2, __A17_1__FO5D, net_U17026_Pad12, TRANmZ, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17027(net_U17026_Pad12, net_R17017_Pad2, net_U17027_Pad3, net_R17018_Pad2, net_U17027_Pad5, net_R17018_Pad2, GND, net_R17018_Pad2, net_U17027_Pad9, CHOR01_n, net_U17027_Pad11, CHOR07_n, net_U17027_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U17028(net_U17026_Pad3, GOJAM, MNIMpR, MNIMmR, TRST9, net_U17027_Pad5, GND, net_U17027_Pad9, TRST10, PCHGOF, ROLGOF, net_U17028_Pad12, __A17_1__TRP31B, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17029(net_U17026_Pad3, net_U17025_Pad10, net_U17028_Pad12, CH3201, MNIMpP, __A17_1__RCH32_n, GND, MNIMmP, __A17_1__RCH32_n, CH3202, MNIMpY, __A17_1__RCH32_n, CH3203, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17030(CH3204, MNIMmY, __A17_1__RCH32_n, CH3205, MNIMpR, __A17_1__RCH32_n, GND, MNIMmR, __A17_1__RCH32_n, CH3206, TRST9, __A17_1__RCH32_n, CH3207, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U17031(CH3208, TRST10, __A17_1__RCH32_n, CH3209, PCHGOF, __A17_1__RCH32_n, GND, ROLGOF, __A17_1__RCH32_n, CH3210, net_U17031_Pad11, net_U17031_Pad12, net_U17031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U17032(net_U17027_Pad3, MNIMpP, MNIMmP, MNIMpY, MNIMmY,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17033(WCHG_n, XT1_n, net_U17033_Pad3, net_R17018_Pad2, F05A_n, net_U17031_Pad11, GND, net_U17031_Pad12, net_U17031_Pad13, __A17_1__FO5D, net_R17018_Pad2, net_U17033_Pad12, XB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U17034(__A17_1__TRP32, net_U17031_Pad13, F05B_n, net_U17034_Pad4, CHWL14_n, WCH13_n, GND, net_U17034_Pad4, net_U17034_Pad9, net_U17033_Pad3, net_U17034_Pad11, TPOR_n, HNDRPT, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17035(net_U17033_Pad3, GOJAM, __A17_1__TRP31A, __A17_1__TRP31B, __A17_1__TRP32, net_U17034_Pad11, GND, net_U17027_Pad11, CH1301, net_U17035_Pad10, CH1401, net_U17034_Pad9, __A17_1__TRP32, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17036(CH3313, PIPAFL, RCH33_n, CH3314, AGCWAR, RCH33_n, GND, OSCALM, RCH33_n, CH3316, CHWL01_n, __A17_2__WCH10_n, net_U17036_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17037(net_U17002_Pad13, net_U17036_Pad13, net_U17037_Pad3, net_U17037_Pad3, net_U17002_Pad13, __A17_2__CCH10, GND, net_U17002_Pad13, __A17_2__RCH10_n, net_U17035_Pad10, CHWL02_n, __A17_2__WCH10_n, net_U17037_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17038(net_U17038_Pad1, net_U17037_Pad13, net_U17038_Pad3, net_U17038_Pad3, net_U17038_Pad1, __A17_2__CCH10, GND, net_U17038_Pad1, __A17_2__RCH10_n, net_U17038_Pad10, CHWL03_n, __A17_2__WCH10_n, net_U17038_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17039(net_U17038_Pad1, RLYB02, net_U17039_Pad3, RLYB03, net_U17039_Pad5, RLYB04, GND, RLYB05, net_U17039_Pad9, RLYB06, net_U17039_Pad11, RLYB07, net_U17039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17040(CH1302, net_U17038_Pad10, CH1303, net_U17040_Pad4, CH1403, net_U17040_Pad6, GND, net_U17040_Pad8, CH1304, net_U17040_Pad10, CH1404, net_U17040_Pad12, CH1402, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17041(net_U17040_Pad12, CHOR02_n, net_U17040_Pad6, CHOR03_n, net_U17040_Pad8, CHOR04_n, GND, CHOR05_n, net_U17041_Pad9, CHOR06_n, net_U17041_Pad11, CHOR08_n, net_U17041_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17042(net_U17039_Pad3, net_U17038_Pad13, net_U17042_Pad3, net_U17042_Pad3, net_U17039_Pad3, __A17_2__CCH10, GND, net_U17039_Pad3, __A17_2__RCH10_n, net_U17040_Pad4, CHWL04_n, __A17_2__WCH10_n, net_U17042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17043(net_U17039_Pad5, net_U17042_Pad13, net_U17043_Pad3, net_U17043_Pad3, net_U17039_Pad5, __A17_2__CCH10, GND, net_U17039_Pad5, __A17_2__RCH10_n, net_U17040_Pad10, CHWL05_n, __A17_2__WCH10_n, net_U17043_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17044(net_U17039_Pad9, net_U17043_Pad13, net_U17044_Pad3, net_U17044_Pad3, net_U17039_Pad9, __A17_2__CCH10, GND, net_U17039_Pad9, __A17_2__RCH10_n, net_U17044_Pad10, CHWL06_n, __A17_2__WCH10_n, net_U17044_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17045(CH1305, net_U17044_Pad10, CH1306, net_U17045_Pad4, CH1406, net_U17041_Pad11, GND,  ,  ,  ,  , net_U17041_Pad9, CH1405, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17046(net_U17039_Pad11, net_U17044_Pad13, net_U17046_Pad3, net_U17046_Pad3, net_U17039_Pad11, __A17_2__CCH10, GND, net_U17039_Pad11, __A17_2__RCH10_n, net_U17045_Pad4, CHWL07_n, __A17_2__WCH10_n, net_U17046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17047(net_U17039_Pad13, net_U17046_Pad13, net_U17047_Pad3, net_U17047_Pad3, net_U17039_Pad13, __A17_2__CCH10, GND, net_U17039_Pad13, __A17_2__RCH10_n, net_U17047_Pad10, CHWL08_n, __A17_2__WCH10_n, net_U17047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17048(CH1307, net_U17047_Pad10, CH1308, net_U17048_Pad4, CH1408, net_U17041_Pad13, GND, net_U17048_Pad8, CH1309, net_U17048_Pad10, CH1409, net_U17027_Pad13, CH1407, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17049(net_U17049_Pad1, net_U17047_Pad13, net_U17049_Pad3, net_U17049_Pad3, net_U17049_Pad1, __A17_2__CCH10, GND, net_U17049_Pad1, __A17_2__RCH10_n, net_U17048_Pad4, CHWL09_n, __A17_2__WCH10_n, net_U17049_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17050(net_U17049_Pad1, RLYB08, net_U17050_Pad3, RLYB09, net_U17050_Pad5, RLYB10, GND, RLYB11, net_U17050_Pad9, RYWD12, net_U17050_Pad11, RYWD13, net_U17050_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17051(net_U17050_Pad3, net_U17049_Pad13, net_U17051_Pad3, net_U17051_Pad3, net_U17050_Pad3, __A17_2__CCH10, GND, net_U17050_Pad3, __A17_2__RCH10_n, net_U17048_Pad10, CHWL10_n, __A17_2__WCH10_n, net_U17051_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17052(net_U17048_Pad8, CHOR09_n, net_U17052_Pad3, CHOR10_n, net_U17052_Pad5, CHOR11_n, GND, CHOR12_n, net_U17052_Pad9, CHOR13_n, net_U17052_Pad11, CHOR14_n, net_U17052_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17053(net_U17050_Pad5, net_U17051_Pad13, net_U17053_Pad3, net_U17053_Pad3, net_U17050_Pad5, __A17_2__CCH10, GND, net_U17050_Pad5, __A17_2__RCH10_n, net_U17053_Pad10, CHWL11_n, __A17_2__WCH10_n, net_U17053_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17054(CH1310, net_U17053_Pad10, CH1311, net_U17054_Pad4, CH1411, net_U17052_Pad5, GND, net_U17052_Pad9, CH3312, net_U17054_Pad10, CH1412, net_U17052_Pad3, CH1410, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17055(net_U17050_Pad9, net_U17053_Pad13, net_U17055_Pad3, net_U17055_Pad3, net_U17050_Pad9, __A17_2__CCH10, GND, net_U17050_Pad9, __A17_2__RCH10_n, net_U17054_Pad4, CHWL12_n, __A17_2__WCH10_n, net_U17055_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17056(net_U17050_Pad11, net_U17055_Pad13, net_U17056_Pad3, net_U17056_Pad3, net_U17050_Pad11, __A17_2__CCH10, GND, net_U17050_Pad11, __A17_2__RCH10_n, net_U17054_Pad10, CHWL13_n, __A17_2__WCH10_n, net_U17056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17057(net_U17050_Pad13, net_U17056_Pad13, net_U17057_Pad3, net_U17057_Pad3, net_U17050_Pad13, __A17_2__CCH10, GND, net_U17050_Pad13, __A17_2__RCH10_n, net_U17057_Pad10, CHWL14_n, __A17_2__WCH10_n, net_U17057_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17058(net_U17058_Pad1, net_U17057_Pad13, net_U17058_Pad3, net_U17058_Pad3, net_U17058_Pad1, __A17_2__CCH10, GND, net_U17058_Pad1, __A17_2__RCH10_n, net_U17058_Pad10, CHWL16_n, __A17_2__WCH10_n, net_U17058_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17059(net_U17058_Pad1, RYWD14, net_U17059_Pad3, RYWD16, net_U17059_Pad5, __A17_2__WCH10_n, GND, __A17_2__CCH10, net_U17059_Pad9, WCH11_n, net_U17033_Pad12, CCH11, net_U17059_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17060(net_U17059_Pad3, net_U17058_Pad13, net_U17060_Pad3, net_U17060_Pad3, net_U17059_Pad3, __A17_2__CCH10, GND, net_U17059_Pad3, __A17_2__RCH10_n, net_U17060_Pad10, net_U17060_Pad11, GOJAM, net_U17059_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17061(net_U17061_Pad1, CHOR16_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2
    U74HC27 U17062(CH1213, net_U17057_Pad10, CH1214, net_U17058_Pad10, CH1414, net_U17052_Pad13, GND, net_U17061_Pad1, CH1316, net_U17060_Pad10, CH1416, net_U17052_Pad11, CH1413, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17063(WCHG_n, XB0_n, CCHG_n, XT1_n, XB0_n, net_U17060_Pad11, GND, net_U17063_Pad8, CCHG_n, XT1_n, XB1_n, net_U17059_Pad5, XT1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17064(net_U17064_Pad1, XT1_n, XB0_n, net_U17059_Pad13, net_U17063_Pad8, GOJAM, GND, XT1_n, XB1_n, net_U17064_Pad10,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17065(net_U17064_Pad1, __A17_2__RCH10_n, net_U17064_Pad10, RCH11_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule