`timescale 1ns/1ps
`default_nettype none

module inout_iii(SIM_RST, SIM_CLK, p4VDC, p4VSW, GND, GOJAM, STOP, T05, T11, F08B, FS09_n, F09A, F09B, F09B_n, F10A, F10A_n, F17A, F17B, SB0_n, SB2_n, F5ASB2_n, F5BSB2_n, CCH13, RCH13_n, WCH13_n, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL11_n, GTSET_n, GTRST_n, MKEY1, MKEY2, MKEY3, MKEY4, MKEY5, MAINRS, NKEY1, NKEY2, NKEY3, NKEY4, NKEY5, NAVRST, MARK, MRKREJ, MRKRST, SBYBUT, LRIN0, LRIN1, RRIN0, RRIN1, XT1_n, XB5_n, XB6_n, ALTEST, TPOR_n, SBY, STNDBY_n, SBYLIT, SBYREL_n, KYRPT1, KYRPT2, MKRPT, RADRPT, RNRADP, RNRADM, CH1301, CH1302, CH1303, CH1304, CH1311, CH1501, CH1502, CH1503, CH1504, CH1505, CH1601, CH1602, CH1603, CH1604, CH1605, CH1606, CH1607);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VDC;
    input wire p4VSW;
    input wire GND;
    input wire ALTEST;
    input wire CCH13;
    output wire CH1301;
    output wire CH1302;
    output wire CH1303;
    output wire CH1304;
    output wire CH1311;
    output wire CH1501;
    output wire CH1502;
    output wire CH1503;
    output wire CH1504;
    output wire CH1505;
    output wire CH1601;
    output wire CH1602;
    output wire CH1603;
    output wire CH1604;
    output wire CH1605;
    output wire CH1606;
    output wire CH1607;
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL11_n;
    input wire F08B;
    input wire F09A;
    input wire F09B;
    input wire F09B_n;
    input wire F10A;
    input wire F10A_n;
    input wire F17A;
    input wire F17B;
    input wire F5ASB2_n;
    input wire F5BSB2_n;
    input wire FS09_n;
    input wire GOJAM;
    input wire GTRST_n;
    input wire GTSET_n;
    output wire KYRPT1;
    output wire KYRPT2;
    input wire LRIN0;
    input wire LRIN1;
    input wire MAINRS;
    input wire MARK;
    input wire MKEY1;
    input wire MKEY2;
    input wire MKEY3;
    input wire MKEY4;
    input wire MKEY5;
    output wire MKRPT;
    input wire MRKREJ;
    input wire MRKRST;
    input wire NAVRST;
    input wire NKEY1;
    input wire NKEY2;
    input wire NKEY3;
    input wire NKEY4;
    input wire NKEY5;
    output wire RADRPT;
    input wire RCH13_n;
    output wire RNRADM;
    output wire RNRADP;
    input wire RRIN0;
    input wire RRIN1;
    input wire SB0_n;
    input wire SB2_n;
    output wire SBY;
    input wire SBYBUT;
    output wire SBYLIT;
    output wire SBYREL_n;
    output wire STNDBY_n;
    input wire STOP;
    input wire T05;
    input wire T11;
    output wire TPOR_n;
    input wire WCH13_n;
    input wire XB5_n;
    input wire XB6_n;
    input wire XT1_n;
    wire __A18_1__F08B_n;
    wire __A18_1__F09A_n;
    wire __A18_1__F09D;
    wire __A18_1__F17A_n;
    wire __A18_1__F17B_n;
    wire __A18_1__RCH15_n;
    wire __A18_1__RCH16_n;
    wire __A18_1__STNDBY;
    wire __A18_2__ACTV_n;
    wire __A18_2__ADVCNT;
    wire __A18_2__CNTOF9; //FPGA#wand
    wire __A18_2__F10AS0;
    wire __A18_2__HERB;
    wire __A18_2__LRRANG;
    wire __A18_2__LRSYNC;
    wire __A18_2__LRXVEL;
    wire __A18_2__LRYVEL;
    wire __A18_2__LRZVEL;
    wire __A18_2__RRRANG;
    wire __A18_2__RRRARA;
    wire __A18_2__RRSYNC;
    wire net_R18001_Pad2; //FPGA#wand
    wire net_R18002_Pad2; //FPGA#wand
    wire net_U18001_Pad1;
    wire net_U18001_Pad12;
    wire net_U18001_Pad13;
    wire net_U18001_Pad3;
    wire net_U18001_Pad6;
    wire net_U18002_Pad10;
    wire net_U18002_Pad11;
    wire net_U18002_Pad12;
    wire net_U18002_Pad2;
    wire net_U18002_Pad4;
    wire net_U18002_Pad5;
    wire net_U18002_Pad6;
    wire net_U18002_Pad8;
    wire net_U18002_Pad9;
    wire net_U18003_Pad13;
    wire net_U18004_Pad10;
    wire net_U18005_Pad13;
    wire net_U18005_Pad3;
    wire net_U18006_Pad10;
    wire net_U18006_Pad12;
    wire net_U18006_Pad6;
    wire net_U18007_Pad11;
    wire net_U18007_Pad13;
    wire net_U18007_Pad5;
    wire net_U18007_Pad9;
    wire net_U18008_Pad10;
    wire net_U18008_Pad11;
    wire net_U18008_Pad13;
    wire net_U18008_Pad3;
    wire net_U18008_Pad6;
    wire net_U18009_Pad2;
    wire net_U18009_Pad3;
    wire net_U18009_Pad8;
    wire net_U18010_Pad12;
    wire net_U18010_Pad13;
    wire net_U18010_Pad5;
    wire net_U18011_Pad1;
    wire net_U18011_Pad10;
    wire net_U18012_Pad1;
    wire net_U18012_Pad12;
    wire net_U18012_Pad13;
    wire net_U18012_Pad3;
    wire net_U18013_Pad10;
    wire net_U18013_Pad11;
    wire net_U18013_Pad12;
    wire net_U18013_Pad2;
    wire net_U18013_Pad4;
    wire net_U18013_Pad5;
    wire net_U18013_Pad6;
    wire net_U18013_Pad8;
    wire net_U18013_Pad9;
    wire net_U18014_Pad13;
    wire net_U18015_Pad10;
    wire net_U18016_Pad3;
    wire net_U18017_Pad10;
    wire net_U18017_Pad6;
    wire net_U18018_Pad13;
    wire net_U18018_Pad4;
    wire net_U18023_Pad10;
    wire net_U18023_Pad6;
    wire net_U18025_Pad10;
    wire net_U18025_Pad11;
    wire net_U18025_Pad2;
    wire net_U18025_Pad4;
    wire net_U18025_Pad5;
    wire net_U18025_Pad6;
    wire net_U18025_Pad8;
    wire net_U18025_Pad9;
    wire net_U18026_Pad13;
    wire net_U18026_Pad3;
    wire net_U18027_Pad11;
    wire net_U18027_Pad12;
    wire net_U18027_Pad13;
    wire net_U18028_Pad12;
    wire net_U18028_Pad13;
    wire net_U18028_Pad5;
    wire net_U18028_Pad9;
    wire net_U18029_Pad10;
    wire net_U18029_Pad11;
    wire net_U18029_Pad8;
    wire net_U18029_Pad9;
    wire net_U18030_Pad1;
    wire net_U18030_Pad10;
    wire net_U18030_Pad11;
    wire net_U18031_Pad10;
    wire net_U18031_Pad11;
    wire net_U18031_Pad12;
    wire net_U18031_Pad3;
    wire net_U18031_Pad4;
    wire net_U18031_Pad5;
    wire net_U18031_Pad8;
    wire net_U18031_Pad9;
    wire net_U18032_Pad1;
    wire net_U18032_Pad13;
    wire net_U18033_Pad13;
    wire net_U18034_Pad1;
    wire net_U18034_Pad13;
    wire net_U18034_Pad3;
    wire net_U18035_Pad1;
    wire net_U18035_Pad3;
    wire net_U18036_Pad10;
    wire net_U18036_Pad12;
    wire net_U18036_Pad13;
    wire net_U18036_Pad3;
    wire net_U18037_Pad11;
    wire net_U18037_Pad8;
    wire net_U18037_Pad9;
    wire net_U18038_Pad12;
    wire net_U18038_Pad13;
    wire net_U18038_Pad4;
    wire net_U18039_Pad12;
    wire net_U18039_Pad13;
    wire net_U18039_Pad9;
    wire net_U18040_Pad10;
    wire net_U18040_Pad12;
    wire net_U18040_Pad13;
    wire net_U18041_Pad3;
    wire net_U18041_Pad5;
    wire net_U18041_Pad6;
    wire net_U18042_Pad12;
    wire net_U18042_Pad13;
    wire net_U18042_Pad4;
    wire net_U18044_Pad10;
    wire net_U18044_Pad13;
    wire net_U18044_Pad9;
    wire net_U18048_Pad1;
    wire net_U18048_Pad10;
    wire net_U18048_Pad12;
    wire net_U18048_Pad13;
    wire net_U18048_Pad4;
    wire net_U18048_Pad6;
    wire net_U18049_Pad9;
    wire net_U18050_Pad10;
    wire net_U18050_Pad12;
    wire net_U18050_Pad5;
    wire net_U18050_Pad8;
    wire net_U18051_Pad10;
    wire net_U18051_Pad4;
    wire net_U18051_Pad5;
    wire net_U18051_Pad6;
    wire net_U18051_Pad8;
    wire net_U18119_Pad1;
    wire net_U18119_Pad10;
    wire net_U18119_Pad11;
    wire net_U18120_Pad13;
    wire net_U18120_Pad2;
    wire net_U18121_Pad1;
    wire net_U18121_Pad10;
    wire net_U18121_Pad12;
    wire net_U18121_Pad13;
    wire net_U18122_Pad1;
    wire net_U18122_Pad10;
    wire net_U18122_Pad13;
    wire net_U18122_Pad3;
    wire net_U18122_Pad8;
    wire net_U18124_Pad1;
    wire net_U18124_Pad4;

    pullup R18001(net_R18001_Pad2);
    pullup R18002(net_R18002_Pad2);
    pullup R18003(__A18_2__CNTOF9);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U18001(net_U18001_Pad1, MKEY1, net_U18001_Pad3, net_U18001_Pad3, net_U18001_Pad1, net_U18001_Pad6, GND, net_U18001_Pad1, __A18_1__RCH15_n, CH1501, MKEY2, net_U18001_Pad12, net_U18001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U18002(net_U18001_Pad1, net_U18002_Pad2, net_U18001_Pad13, net_U18002_Pad4, net_U18002_Pad5, net_U18002_Pad6, GND, net_U18002_Pad8, net_U18002_Pad9, net_U18002_Pad10, net_U18002_Pad11, net_U18002_Pad12, MAINRS, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18003(net_U18001_Pad12, net_U18001_Pad13, net_U18001_Pad6, CH1502, net_U18001_Pad13, __A18_1__RCH15_n, GND, MKEY3, net_U18003_Pad13, net_U18002_Pad5, net_U18002_Pad5, net_U18001_Pad6, net_U18003_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18004(CH1503, net_U18002_Pad5, __A18_1__RCH15_n, net_U18002_Pad9, MKEY4, net_U18004_Pad10, GND, net_U18002_Pad9, net_U18001_Pad6, net_U18004_Pad10, net_U18002_Pad9, __A18_1__RCH15_n, CH1504, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18005(net_U18002_Pad11, MKEY5, net_U18005_Pad3, net_U18005_Pad3, net_U18002_Pad11, net_U18001_Pad6, GND, net_U18002_Pad11, __A18_1__RCH15_n, CH1505, net_U18002_Pad8, net_U18002_Pad10, net_U18005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18006(net_U18002_Pad2, net_U18002_Pad4, net_U18006_Pad10, net_R18001_Pad2, __A18_1__F09D, net_U18006_Pad6, GND, KYRPT1, TPOR_n, net_U18006_Pad10, F09B_n, net_U18006_Pad12, net_U18002_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U18007(net_U18006_Pad12, net_R18001_Pad2, net_U18005_Pad13, net_R18001_Pad2, net_U18007_Pad5, net_R18002_Pad2, GND, net_R18002_Pad2, net_U18007_Pad9, __A18_2__CNTOF9, net_U18007_Pad11, __A18_2__CNTOF9, net_U18007_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U18008(net_U18002_Pad12, net_U18001_Pad6, net_U18008_Pad3, __A18_1__RCH15_n, net_R18001_Pad2, net_U18008_Pad6, GND, net_U18008_Pad11, NAVRST, net_U18008_Pad10, net_U18008_Pad11, __A18_1__RCH16_n, net_U18008_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18009(__A18_2__RRSYNC, net_U18009_Pad2, net_U18009_Pad3, net_U18008_Pad3, XT1_n, XB5_n, GND, net_U18009_Pad8, net_U18006_Pad6, net_U18006_Pad10, T05, T11, TPOR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U18010(net_U18009_Pad8, __A18_1__F09A_n, net_R18001_Pad2, net_U18001_Pad6, net_U18010_Pad5,  , GND,  , __A18_1__F09A_n, net_R18002_Pad2, net_U18008_Pad10, net_U18010_Pad12, net_U18010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18011(net_U18011_Pad1, net_U18008_Pad6, net_U18002_Pad12, net_U18010_Pad5, net_U18011_Pad1, net_U18011_Pad10, GND, net_U18010_Pad5, KYRPT1, net_U18011_Pad10, XT1_n, XB6_n, net_U18008_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U18012(net_U18012_Pad1, NKEY1, net_U18012_Pad3, net_U18012_Pad3, net_U18012_Pad1, net_U18008_Pad10, GND, net_U18012_Pad1, __A18_1__RCH16_n, CH1601, NKEY2, net_U18012_Pad12, net_U18012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U18013(net_U18012_Pad1, net_U18013_Pad2, net_U18012_Pad13, net_U18013_Pad4, net_U18013_Pad5, net_U18013_Pad6, GND, net_U18013_Pad8, net_U18013_Pad9, net_U18013_Pad10, net_U18013_Pad11, net_U18013_Pad12, net_R18002_Pad2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18014(net_U18012_Pad12, net_U18012_Pad13, net_U18008_Pad10, CH1602, net_U18012_Pad13, __A18_1__RCH16_n, GND, NKEY3, net_U18014_Pad13, net_U18013_Pad5, net_U18013_Pad5, net_U18008_Pad10, net_U18014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18015(CH1603, net_U18013_Pad5, __A18_1__RCH16_n, net_U18013_Pad9, NKEY4, net_U18015_Pad10, GND, net_U18013_Pad9, net_U18008_Pad10, net_U18015_Pad10, net_U18013_Pad9, __A18_1__RCH16_n, CH1604, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18016(net_U18013_Pad11, NKEY5, net_U18016_Pad3, net_U18016_Pad3, net_U18013_Pad11, net_U18008_Pad10, GND, net_U18013_Pad11, __A18_1__RCH16_n, CH1605, net_U18013_Pad8, net_U18013_Pad10, net_U18007_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18017(net_U18013_Pad2, net_U18013_Pad4, net_U18017_Pad10, net_R18002_Pad2, __A18_1__F09D, net_U18017_Pad6, GND, KYRPT2, TPOR_n, net_U18017_Pad10, F09B_n, net_U18007_Pad5, net_U18013_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18018(net_U18017_Pad10, net_U18010_Pad13, net_U18017_Pad6, net_U18018_Pad4, net_U18013_Pad12, net_U18008_Pad11, GND, net_U18018_Pad4, net_U18018_Pad13, net_U18010_Pad12, net_U18010_Pad12, KYRPT2, net_U18018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18119(net_U18119_Pad1, WCH13_n, CHWL11_n, net_U18119_Pad11, net_U18119_Pad1, net_U18119_Pad10, GND, net_U18119_Pad11, CCH13, net_U18119_Pad10, net_U18119_Pad11, RCH13_n, CH1311, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U18120(SBYBUT, net_U18120_Pad2, F17A, __A18_1__F17A_n, F17B, __A18_1__F17B_n, GND, STNDBY_n, __A18_1__STNDBY, SBY, STNDBY_n, SBYLIT, net_U18120_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18121(net_U18121_Pad1, __A18_1__F17A_n, net_U18120_Pad2, net_U18121_Pad12, net_U18121_Pad1, net_U18121_Pad10, GND, net_U18121_Pad12, net_U18120_Pad2, net_U18121_Pad10, __A18_1__F17B_n, net_U18121_Pad12, net_U18121_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18122(net_U18122_Pad1, net_U18121_Pad13, net_U18122_Pad3, net_U18122_Pad3, net_U18122_Pad1, net_U18120_Pad2, GND, net_U18122_Pad8, net_U18122_Pad13, net_U18122_Pad10, net_U18122_Pad10, net_U18122_Pad1, net_U18122_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U18023( ,  , __A18_2__ACTV_n, RADRPT, CCH13, net_U18023_Pad6, GND, __A18_2__ADVCNT, F10A_n, net_U18023_Pad10, SB2_n,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18124(net_U18124_Pad1, net_U18122_Pad13, net_U18122_Pad1, net_U18124_Pad4, net_U18122_Pad13, __A18_1__STNDBY, GND, net_U18124_Pad4, net_U18124_Pad1, __A18_1__STNDBY, __A18_1__STNDBY, ALTEST, net_U18120_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U18025(MRKRST, net_U18025_Pad2, net_U18025_Pad2, net_U18025_Pad4, net_U18025_Pad5, net_U18025_Pad6, GND, net_U18025_Pad8, net_U18025_Pad9, net_U18025_Pad10, net_U18025_Pad11, __A18_1__F08B_n, F08B, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18026(net_U18025_Pad5, MARK, net_U18026_Pad3, net_U18026_Pad3, net_U18025_Pad5, net_U18025_Pad4, GND, MRKREJ, net_U18026_Pad13, net_U18025_Pad9, net_U18025_Pad9, net_U18025_Pad4, net_U18026_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U18027(CH1606, net_U18025_Pad5, __A18_1__RCH16_n, CH1607, net_U18025_Pad9, __A18_1__RCH16_n, GND, net_U18025_Pad6, net_U18025_Pad8, net_U18025_Pad11, net_U18027_Pad11, net_U18027_Pad12, net_U18027_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U18028(net_U18027_Pad11, __A18_1__F09A_n, net_U18025_Pad11, net_U18025_Pad4, net_U18028_Pad5,  , GND,  , net_U18028_Pad9, RADRPT, __A18_2__ADVCNT, net_U18028_Pad12, net_U18028_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18029(TPOR_n, net_U18027_Pad13, net_U18027_Pad13, net_U18025_Pad11, __A18_1__F09D, net_U18027_Pad12, GND, net_U18029_Pad8, net_U18029_Pad9, net_U18029_Pad10, net_U18029_Pad11, MKRPT, F09B_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18030(net_U18030_Pad1, net_U18025_Pad10, net_U18025_Pad2, net_U18028_Pad5, net_U18030_Pad1, net_U18030_Pad10, GND, net_U18028_Pad5, MKRPT, net_U18030_Pad10, net_U18030_Pad11, FS09_n, __A18_1__F09D, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1) U18031(__A18_1__F08B_n, net_U18030_Pad11, net_U18031_Pad3, net_U18031_Pad4, net_U18031_Pad5, net_U18029_Pad9, GND, net_U18031_Pad8, net_U18031_Pad9, net_U18031_Pad10, net_U18031_Pad11, net_U18031_Pad12, __A18_2__CNTOF9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18032(net_U18032_Pad1, CHWL04_n, WCH13_n, __A18_2__ACTV_n, net_U18032_Pad1, net_U18023_Pad6, GND, RCH13_n, __A18_2__ACTV_n, CH1304, CHWL03_n, WCH13_n, net_U18032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18033(net_U18031_Pad3, net_U18032_Pad13, net_U18031_Pad5, net_U18031_Pad5, net_U18031_Pad3, CCH13, GND, RCH13_n, net_U18031_Pad3, CH1303, CHWL02_n, WCH13_n, net_U18033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18034(net_U18034_Pad1, net_U18033_Pad13, net_U18034_Pad3, net_U18034_Pad3, net_U18034_Pad1, CCH13, GND, RCH13_n, net_U18034_Pad1, CH1302, CHWL01_n, WCH13_n, net_U18034_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18035(net_U18035_Pad1, net_U18034_Pad13, net_U18035_Pad3, net_U18035_Pad3, net_U18035_Pad1, CCH13, GND, RCH13_n, net_U18035_Pad1, CH1301, F10A_n, SB0_n, __A18_2__F10AS0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18036(net_U18023_Pad10, __A18_2__F10AS0, net_U18036_Pad3, net_U18036_Pad3, net_U18023_Pad10, __A18_2__ACTV_n, GND, net_U18028_Pad12, net_U18036_Pad12, net_U18036_Pad10, net_U18028_Pad13, net_U18036_Pad12, net_U18036_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18037(net_U18028_Pad13, __A18_2__ADVCNT, net_U18036_Pad13, RADRPT, net_U18028_Pad13, net_U18028_Pad9, GND, net_U18037_Pad8, net_U18037_Pad9, net_U18028_Pad9, net_U18037_Pad11, net_U18028_Pad12, net_U18036_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18038(net_U18036_Pad12, net_U18036_Pad13, net_U18028_Pad12, net_U18038_Pad4, net_U18038_Pad13, net_U18037_Pad9, GND, net_U18037_Pad8, net_U18038_Pad12, net_U18037_Pad11, net_U18037_Pad9, net_U18038_Pad12, net_U18038_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U18039(net_U18037_Pad9, net_U18038_Pad4, RADRPT, net_U18028_Pad9, net_U18037_Pad8,  , GND,  , net_U18039_Pad9, RADRPT, net_U18038_Pad4, net_U18039_Pad12, net_U18039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18040(net_U18038_Pad12, net_U18038_Pad13, net_U18037_Pad8, net_U18039_Pad9, net_U18040_Pad13, net_U18039_Pad13, GND, net_U18039_Pad12, net_U18040_Pad12, net_U18040_Pad10, net_U18039_Pad13, net_U18040_Pad12, net_U18040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18041(net_U18039_Pad13, net_U18038_Pad4, net_U18041_Pad3, net_U18039_Pad9, net_U18041_Pad5, net_U18041_Pad6, GND, net_U18007_Pad13, net_U18038_Pad12, net_U18036_Pad13, F10A, net_U18039_Pad12, net_U18040_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18042(net_U18040_Pad12, net_U18040_Pad13, net_U18039_Pad12, net_U18042_Pad4, net_U18042_Pad13, net_U18041_Pad3, GND, net_U18041_Pad6, net_U18042_Pad12, net_U18041_Pad5, net_U18041_Pad3, net_U18042_Pad12, net_U18042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U18043(net_U18041_Pad3, net_U18042_Pad4, RADRPT, net_U18039_Pad9, net_U18041_Pad6,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U18044(net_U18042_Pad12, net_U18042_Pad13, net_U18041_Pad6, net_U18007_Pad11, net_U18042_Pad13, net_U18040_Pad12, GND, __A18_2__ADVCNT, net_U18044_Pad9, net_U18044_Pad10, net_U18034_Pad3, net_U18035_Pad3, net_U18044_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18045(net_U18044_Pad10, __A18_2__CNTOF9, net_U18031_Pad4, net_U18044_Pad10, F5BSB2_n, net_U18031_Pad9, GND, net_U18031_Pad11, F5BSB2_n, net_U18044_Pad10, net_U18029_Pad9, net_U18044_Pad9, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18046(net_U18034_Pad3, net_U18035_Pad1, net_U18031_Pad8, net_U18035_Pad3, net_U18034_Pad1, __A18_2__RRRARA, GND, __A18_2__LRXVEL, net_U18035_Pad3, net_U18034_Pad3, net_U18031_Pad10, __A18_2__RRRANG, net_U18031_Pad8, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18047(net_U18031_Pad10, net_U18035_Pad1, net_U18031_Pad10, net_U18034_Pad1, net_U18035_Pad3, __A18_2__LRZVEL, GND, __A18_2__LRRANG, net_U18031_Pad10, net_U18034_Pad1, net_U18035_Pad1, __A18_2__LRYVEL, net_U18034_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U18048(net_U18048_Pad1, net_U18031_Pad12, GTSET_n, net_U18048_Pad4, net_U18048_Pad1, net_U18048_Pad6, GND, F5ASB2_n, net_U18048_Pad4, net_U18048_Pad10, net_U18048_Pad10, net_U18048_Pad12, net_U18048_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18049(net_U18048_Pad4, RADRPT, net_U18048_Pad13, F09B, GOJAM, net_U18048_Pad12, GND, RADRPT, net_U18049_Pad9, net_U18048_Pad13, GTRST_n, net_U18048_Pad6, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U18050(TPOR_n, __A18_2__HERB, __A18_2__HERB, net_U18049_Pad9, net_U18050_Pad5, net_U18009_Pad2, GND, net_U18050_Pad8, RRIN1, net_U18050_Pad10, RRIN0, net_U18050_Pad12, LRIN1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U18051(net_U18050_Pad5, net_U18044_Pad13, net_U18031_Pad4, net_U18051_Pad4, net_U18051_Pad5, net_U18051_Pad6, GND, net_U18051_Pad8, net_U18029_Pad8, net_U18051_Pad10, net_U18009_Pad3, net_U18029_Pad9, __A18_2__LRSYNC, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18052(net_U18009_Pad2, net_U18050_Pad8, net_U18009_Pad2, net_U18050_Pad10, net_U18029_Pad11, net_U18051_Pad8, GND, net_U18051_Pad6, net_U18029_Pad9, net_U18050_Pad12, net_U18029_Pad11, net_U18051_Pad5, net_U18029_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U18053(LRIN0, net_U18029_Pad10, net_U18023_Pad6, net_U18029_Pad11, F09A, __A18_1__F09A_n, GND, RNRADP, net_U18051_Pad4, RNRADM, net_U18051_Pad10, net_U18009_Pad3, net_U18048_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U18154(SBY, SBYREL_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U18155(net_U18122_Pad1, STOP,  ,  ,  ,  , GND,  ,  ,  ,  , net_U18122_Pad8, net_U18119_Pad11, p4VDC, SIM_RST, SIM_CLK);
endmodule