`timescale 1ns/1ps
`default_nettype none

module inout_vi(SIM_RST, SIM_CLK, p4VSW, GND, P04_n, SB2_n, F18A, F18B, F5ASB0_n, F5ASB2, F5ASB2_n, CCHG_n, WCHG_n, CCH11, CCH12, CCH13, CCH14, CCH33, RCH11_n, RCH12_n, RCH13_n, RCH14_n, WCH11_n, WCH12_n, WCH13_n, WCH14_n, POUT_n, MOUT_n, ZOUT_n, T6RPT, PIPPLS_n, PIPAXp, PIPAXm, PIPAYp, PIPAYm, PIPAZp, PIPAZm, OCTAD5, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CHWL16_n, XT0_n, XB0_n, XB1_n, XB2_n, XB3_n, XB4_n, XB7_n, T6ON_n, ALTEST, E5, E6, E7_n, CDUXD, CDUYD, CDUZD, PIPAFL, PIPXP, PIPXM, PIPYP, PIPYM, PIPZP, PIPZM, TRUND, SHAFTD, CH0705, CH0706, CH0707, CH1310, CH1316, CH1411, CH1412, CH1413, CH1414, CH1416, CH1108, CH1113, CH1114, CH1116, CH1216, CDUXDP, CDUXDM, CDUYDP, CDUYDM, CDUZDP, CDUZDM);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    output wire ALTEST;
    input wire CCH11;
    input wire CCH12;
    input wire CCH13;
    input wire CCH14;
    input wire CCH33;
    input wire CCHG_n;
    output wire CDUXD;
    output wire CDUXDM;
    output wire CDUXDP;
    output wire CDUYD;
    output wire CDUYDM;
    output wire CDUYDP;
    output wire CDUZD;
    output wire CDUZDM;
    output wire CDUZDP;
    output wire CH0705;
    output wire CH0706;
    output wire CH0707;
    output wire CH1108;
    output wire CH1113;
    output wire CH1114;
    output wire CH1116;
    output wire CH1216;
    output wire CH1310;
    output wire CH1316;
    output wire CH1411;
    output wire CH1412;
    output wire CH1413;
    output wire CH1414;
    output wire CH1416;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire CHWL16_n;
    output wire E5;
    output wire E6;
    output wire E7_n;
    input wire F18A;
    input wire F18B;
    input wire F5ASB0_n;
    input wire F5ASB2;
    input wire F5ASB2_n;
    input wire MOUT_n;
    input wire OCTAD5;
    input wire P04_n;
    output wire PIPAFL;
    input wire PIPAXm;
    input wire PIPAXp;
    input wire PIPAYm;
    input wire PIPAYp;
    input wire PIPAZm;
    input wire PIPAZp;
    input wire PIPPLS_n;
    output wire PIPXM;
    output wire PIPXP;
    output wire PIPYM;
    output wire PIPYP;
    output wire PIPZM;
    output wire PIPZP;
    input wire POUT_n;
    input wire RCH11_n;
    input wire RCH12_n;
    input wire RCH13_n;
    input wire RCH14_n;
    input wire SB2_n;
    output wire SHAFTD;
    output wire T6ON_n;
    input wire T6RPT;
    output wire TRUND;
    input wire WCH11_n;
    input wire WCH12_n;
    input wire WCH13_n;
    input wire WCH14_n;
    input wire WCHG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    input wire XB4_n;
    input wire XB7_n;
    input wire XT0_n;
    input wire ZOUT_n;
    wire __A23_1__BOTHX;
    wire __A23_1__BOTHY;
    wire __A23_1__BOTHZ;
    wire __A23_1__F18AX;
    wire __A23_1__F18A_n;
    wire __A23_1__F18B_n;
    wire __A23_1__MISSX;
    wire __A23_1__MISSY;
    wire __A23_1__MISSZ;
    wire __A23_1__NOXM;
    wire __A23_1__NOXP;
    wire __A23_1__NOYM;
    wire __A23_1__NOYP;
    wire __A23_1__NOZM;
    wire __A23_1__NOZP;
    wire __A23_1__P04A;
    wire __A23_1__PIPAXm_n;
    wire __A23_1__PIPAXp_n;
    wire __A23_1__PIPAYm_n;
    wire __A23_1__PIPAYp_n;
    wire __A23_1__PIPAZm_n;
    wire __A23_1__PIPAZp_n;
    wire __A23_1__PIPGXm;
    wire __A23_1__PIPGXp;
    wire __A23_1__PIPGYm;
    wire __A23_1__PIPGYp;
    wire __A23_1__PIPGZm;
    wire __A23_1__PIPGZp;
    wire __A23_1__PIPSAM;
    wire __A23_1__PIPSAM_n;
    wire __A23_2__CCH07;
    wire __A23_2__ISSTDC;
    wire __A23_2__OT1108;
    wire __A23_2__OT1113;
    wire __A23_2__OT1114;
    wire __A23_2__OT1116;
    wire __A23_2__RCH07_n;
    wire __A23_2__SHFTDM;
    wire __A23_2__SHFTDP;
    wire __A23_2__TRNDM;
    wire __A23_2__TRNDP;
    wire __A23_2__WCH07_n;
    wire net_R23001_Pad2; //FPGA#wand
    wire net_R23002_Pad2; //FPGA#wand
    wire net_U23001_Pad12;
    wire net_U23001_Pad6;
    wire net_U23001_Pad8;
    wire net_U23002_Pad5;
    wire net_U23002_Pad9;
    wire net_U23003_Pad10;
    wire net_U23003_Pad12;
    wire net_U23003_Pad4;
    wire net_U23003_Pad6;
    wire net_U23003_Pad8;
    wire net_U23004_Pad1;
    wire net_U23004_Pad11;
    wire net_U23004_Pad12;
    wire net_U23004_Pad13;
    wire net_U23004_Pad4;
    wire net_U23005_Pad10;
    wire net_U23005_Pad8;
    wire net_U23005_Pad9;
    wire net_U23006_Pad13;
    wire net_U23007_Pad10;
    wire net_U23007_Pad11;
    wire net_U23008_Pad10;
    wire net_U23008_Pad11;
    wire net_U23008_Pad13;
    wire net_U23008_Pad6;
    wire net_U23008_Pad8;
    wire net_U23009_Pad12;
    wire net_U23009_Pad6;
    wire net_U23009_Pad8;
    wire net_U23010_Pad11;
    wire net_U23011_Pad13;
    wire net_U23012_Pad10;
    wire net_U23012_Pad3;
    wire net_U23014_Pad10;
    wire net_U23014_Pad12;
    wire net_U23014_Pad13;
    wire net_U23014_Pad3;
    wire net_U23014_Pad6;
    wire net_U23014_Pad8;
    wire net_U23015_Pad10;
    wire net_U23015_Pad12;
    wire net_U23015_Pad6;
    wire net_U23015_Pad8;
    wire net_U23016_Pad1;
    wire net_U23016_Pad10;
    wire net_U23016_Pad11;
    wire net_U23016_Pad12;
    wire net_U23016_Pad13;
    wire net_U23017_Pad11;
    wire net_U23017_Pad12;
    wire net_U23017_Pad13;
    wire net_U23018_Pad4;
    wire net_U23018_Pad6;
    wire net_U23018_Pad8;
    wire net_U23019_Pad1;
    wire net_U23019_Pad4;
    wire net_U23020_Pad13;
    wire net_U23021_Pad3;
    wire net_U23022_Pad10;
    wire net_U23022_Pad11;
    wire net_U23022_Pad8;
    wire net_U23023_Pad1;
    wire net_U23023_Pad12;
    wire net_U23023_Pad6;
    wire net_U23023_Pad8;
    wire net_U23024_Pad11;
    wire net_U23024_Pad12;
    wire net_U23024_Pad2;
    wire net_U23024_Pad6;
    wire net_U23025_Pad1;
    wire net_U23025_Pad13;
    wire net_U23025_Pad3;
    wire net_U23026_Pad12;
    wire net_U23026_Pad13;
    wire net_U23027_Pad13;
    wire net_U23027_Pad3;
    wire net_U23028_Pad1;
    wire net_U23028_Pad10;
    wire net_U23028_Pad4;
    wire net_U23029_Pad13;
    wire net_U23030_Pad11;
    wire net_U23030_Pad3;
    wire net_U23030_Pad5;
    wire net_U23030_Pad6;
    wire net_U23030_Pad8;
    wire net_U23030_Pad9;
    wire net_U23031_Pad12;
    wire net_U23031_Pad13;
    wire net_U23032_Pad10;
    wire net_U23032_Pad11;
    wire net_U23032_Pad12;
    wire net_U23032_Pad13;
    wire net_U23032_Pad2;
    wire net_U23032_Pad5;
    wire net_U23032_Pad6;
    wire net_U23032_Pad8;
    wire net_U23032_Pad9;
    wire net_U23033_Pad13;
    wire net_U23035_Pad13;
    wire net_U23036_Pad1;
    wire net_U23036_Pad3;
    wire net_U23037_Pad11;
    wire net_U23037_Pad13;
    wire net_U23037_Pad3;
    wire net_U23037_Pad5;
    wire net_U23037_Pad6;
    wire net_U23037_Pad8;
    wire net_U23037_Pad9;
    wire net_U23038_Pad13;
    wire net_U23040_Pad13;
    wire net_U23042_Pad13;
    wire net_U23043_Pad1;
    wire net_U23043_Pad13;
    wire net_U23044_Pad1;
    wire net_U23044_Pad13;
    wire net_U23045_Pad13;
    wire net_U23045_Pad3;
    wire net_U23046_Pad12;
    wire net_U23046_Pad8;
    wire net_U23047_Pad11;
    wire net_U23047_Pad13;
    wire net_U23047_Pad5;
    wire net_U23047_Pad9;
    wire net_U23048_Pad1;
    wire net_U23048_Pad10;
    wire net_U23049_Pad1;
    wire net_U23049_Pad10;
    wire net_U23050_Pad1;
    wire net_U23050_Pad10;
    wire net_U23051_Pad1;
    wire net_U23051_Pad10;
    wire net_U23052_Pad1;
    wire net_U23052_Pad10;
    wire net_U23052_Pad12;
    wire net_U23053_Pad5;
    wire net_U23054_Pad1;
    wire net_U23054_Pad13;
    wire net_U23055_Pad3;

    pullup R23001(net_R23001_Pad2);
    pullup R23002(net_R23002_Pad2);
    U74HC27 #(1'b1, 1'b1, 1'b1) U23001(__A23_1__NOXP, __A23_1__NOXM, __A23_1__NOYM, __A23_1__NOZP, __A23_1__NOZM, net_U23001_Pad6, GND, net_U23001_Pad8, __A23_1__MISSX, __A23_1__MISSY, __A23_1__MISSZ, net_U23001_Pad12, __A23_1__NOYP, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U23002(net_U23001_Pad12, net_R23001_Pad2, net_U23001_Pad6, net_R23001_Pad2, net_U23002_Pad5, net_R23002_Pad2, GND, net_R23002_Pad2, net_U23002_Pad9,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1) U23003(F18B, __A23_1__F18B_n, __A23_1__PIPGXp, net_U23003_Pad4, __A23_1__PIPGXm, net_U23003_Pad6, GND, net_U23003_Pad8, F5ASB2, net_U23003_Pad10, __A23_1__PIPGYp, net_U23003_Pad12, __A23_1__PIPGYm, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23004(net_U23004_Pad1, __A23_1__F18B_n, net_R23001_Pad2, net_U23004_Pad4, F5ASB0_n, net_U23001_Pad8, GND, net_R23002_Pad2, CCH33, PIPAFL, net_U23004_Pad11, net_U23004_Pad12, net_U23004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U23005(__A23_1__BOTHX, __A23_1__BOTHY, net_U23004_Pad1, net_U23004_Pad4, PIPAFL, net_U23002_Pad9, GND, net_U23005_Pad8, net_U23005_Pad9, net_U23005_Pad10, net_U23003_Pad4, net_U23002_Pad5, __A23_1__BOTHZ, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23006(net_U23003_Pad6, net_U23005_Pad10, PIPPLS_n, SB2_n, __A23_1__P04A, __A23_1__PIPSAM, GND,  ,  ,  ,  , net_U23004_Pad11, net_U23006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23007(net_U23004_Pad12, net_U23004_Pad13, net_U23005_Pad8, net_U23007_Pad11, net_U23003_Pad8, net_U23004_Pad13, GND, net_U23004_Pad12, net_U23003_Pad8, net_U23007_Pad10, net_U23007_Pad11, net_U23006_Pad13, net_U23005_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23008(net_U23006_Pad13, net_U23005_Pad9, net_U23007_Pad10, net_U23008_Pad11, net_U23003_Pad8, net_U23008_Pad6, GND, net_U23008_Pad8, net_U23003_Pad8, net_U23008_Pad10, net_U23008_Pad11, net_U23005_Pad10, net_U23008_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23009(net_U23006_Pad13, net_U23005_Pad10, net_U23005_Pad9, net_U23005_Pad10, net_U23003_Pad6, net_U23009_Pad6, GND, net_U23009_Pad8, net_U23006_Pad13, net_U23008_Pad13, net_U23003_Pad6, net_U23009_Pad12, net_U23003_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U23010(net_U23005_Pad9, net_U23008_Pad13, net_U23009_Pad12, net_U23009_Pad6, net_U23008_Pad8, net_U23008_Pad6, GND, net_U23008_Pad8, net_U23008_Pad6, net_U23009_Pad8, net_U23010_Pad11, net_U23010_Pad11, net_U23003_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U23011(net_U23005_Pad10, net_U23008_Pad13, net_U23008_Pad10, __A23_1__BOTHX, net_U23003_Pad6, net_U23003_Pad4, GND, __A23_1__PIPGXm, net_U23011_Pad13, __A23_1__NOXM, __A23_1__NOXM, __A23_1__F18AX, net_U23011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23012(__A23_1__NOXP, __A23_1__PIPGXp, net_U23012_Pad3, net_U23012_Pad3, __A23_1__NOXP, __A23_1__F18AX, GND, __A23_1__MISSX, F5ASB2, net_U23012_Pad10, net_U23003_Pad12, net_U23003_Pad10, __A23_1__BOTHY, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U23013(__A23_1__PIPGXp, __A23_1__PIPGXm, net_U23006_Pad13, net_U23008_Pad13, net_U23003_Pad4, PIPXP, GND, PIPXM, net_U23005_Pad9, net_U23008_Pad13, net_U23003_Pad6, __A23_1__MISSX, net_U23012_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23014(net_U23003_Pad12, net_U23014_Pad10, net_U23014_Pad3, net_U23014_Pad10, net_U23003_Pad10, net_U23014_Pad6, GND, net_U23014_Pad8, net_U23014_Pad13, net_U23014_Pad10, net_U23003_Pad10, net_U23014_Pad12, net_U23014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23015(net_U23014_Pad3, net_U23014_Pad10, net_U23014_Pad13, net_U23015_Pad10, net_U23003_Pad12, net_U23015_Pad6, GND, net_U23015_Pad8, net_U23014_Pad3, net_U23015_Pad10, net_U23003_Pad10, net_U23015_Pad12, net_U23003_Pad12, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23016(net_U23016_Pad1, net_U23014_Pad12, net_U23016_Pad11, net_U23016_Pad11, net_U23016_Pad1, net_U23014_Pad6, GND, net_U23016_Pad12, net_U23016_Pad1, net_U23016_Pad10, net_U23016_Pad11, net_U23016_Pad12, net_U23016_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U23017(net_U23014_Pad8, net_U23015_Pad12, net_U23017_Pad12, net_U23015_Pad6, net_U23015_Pad8, net_U23017_Pad13, GND, __A23_1__MISSY, __A23_1__PIPGYp, __A23_1__PIPGYm, net_U23017_Pad11, net_U23017_Pad12, net_U23017_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U23018(F5ASB2, net_U23016_Pad12, __A23_1__PIPGZp, net_U23018_Pad4, __A23_1__PIPGZm, net_U23018_Pad6, GND, net_U23018_Pad8, F5ASB2, __A23_1__F18A_n, F18A, __A23_1__F18AX, __A23_1__F18A_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U23019(net_U23019_Pad1, net_U23016_Pad12, net_U23017_Pad12, net_U23019_Pad4, net_U23017_Pad13, net_U23016_Pad12, GND, net_U23016_Pad10, net_U23014_Pad13, net_U23014_Pad3, net_U23014_Pad3, net_U23016_Pad13, net_U23014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U23020(net_U23015_Pad10, net_U23019_Pad1, net_U23014_Pad10, net_U23014_Pad10, net_U23015_Pad10, net_U23019_Pad4, GND, __A23_1__PIPGYm, net_U23020_Pad13, __A23_1__NOYM, __A23_1__NOYM, __A23_1__F18AX, net_U23020_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23021(__A23_1__NOYP, __A23_1__PIPGYp, net_U23021_Pad3, net_U23021_Pad3, __A23_1__NOYP, __A23_1__F18AX, GND, __A23_1__MISSY, F5ASB2, net_U23017_Pad11, net_U23018_Pad6, net_U23018_Pad4, __A23_1__BOTHZ, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23022(net_U23014_Pad13, net_U23015_Pad10, net_U23014_Pad3, net_U23015_Pad10, net_U23003_Pad12, PIPYM, GND, net_U23022_Pad8, net_U23018_Pad6, net_U23022_Pad10, net_U23022_Pad11, PIPYP, net_U23003_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23023(net_U23023_Pad1, net_U23022_Pad10, net_U23022_Pad11, net_U23022_Pad10, net_U23018_Pad4, net_U23023_Pad6, GND, net_U23023_Pad8, net_U23023_Pad1, net_U23022_Pad10, net_U23018_Pad6, net_U23023_Pad12, net_U23018_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U23024(net_U23022_Pad11, net_U23024_Pad2, net_U23023_Pad1, net_U23024_Pad2, net_U23018_Pad4, net_U23024_Pad6, GND, __A23_1__MISSZ, __A23_1__PIPGZp, __A23_1__PIPGZm, net_U23024_Pad11, net_U23024_Pad12, net_U23018_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U23025(net_U23025_Pad1, net_U23022_Pad8, net_U23025_Pad3, net_U23025_Pad3, net_U23025_Pad1, net_U23023_Pad12, GND, __A23_1__PIPGZm, net_U23025_Pad13, __A23_1__NOZM, __A23_1__NOZM, __A23_1__F18AX, net_U23025_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U23026(net_U23023_Pad6, net_U23023_Pad8, net_U23026_Pad12, net_U23024_Pad12, net_U23024_Pad6, net_U23026_Pad13, GND, PIPZP, net_U23022_Pad11, net_U23024_Pad2, net_U23018_Pad4, net_U23026_Pad12, net_U23026_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23027(__A23_1__NOZP, __A23_1__PIPGZp, net_U23027_Pad3, net_U23027_Pad3, __A23_1__NOZP, __A23_1__F18AX, GND, __A23_1__MISSZ, F5ASB2, net_U23024_Pad11, net_U23018_Pad8, net_U23025_Pad1, net_U23027_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23028(net_U23028_Pad1, net_U23025_Pad3, net_U23018_Pad8, net_U23028_Pad4, net_U23018_Pad8, net_U23026_Pad12, GND, net_U23026_Pad13, net_U23018_Pad8, net_U23028_Pad10, net_U23027_Pad13, net_U23022_Pad11, net_U23023_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U23029(net_U23022_Pad11, net_U23023_Pad1, net_U23028_Pad1, net_U23024_Pad2, net_U23028_Pad4, net_U23022_Pad10, GND, net_U23024_Pad2, net_U23028_Pad10, net_U23022_Pad10, CHWL16_n, WCH14_n, net_U23029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23030(net_U23023_Pad1, net_U23024_Pad2, net_U23030_Pad3, CCH14, net_U23030_Pad5, net_U23030_Pad6, GND, net_U23030_Pad8, net_U23030_Pad9, CCH14, net_U23030_Pad11, PIPZM, net_U23018_Pad6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23031(net_U23030_Pad3, net_U23029_Pad13, net_U23030_Pad6, CH1416, RCH14_n, net_U23030_Pad3, GND, net_U23030_Pad3, F5ASB2_n, CDUXD, XB0_n, net_U23031_Pad12, net_U23031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0) U23032(net_U23031_Pad13, net_U23032_Pad2, OCTAD5, net_U23031_Pad12, net_U23032_Pad5, net_U23032_Pad6, GND, net_U23032_Pad8, net_U23032_Pad9, net_U23032_Pad10, net_U23032_Pad11, net_U23032_Pad12, net_U23032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23033(CDUXDP, POUT_n, net_U23032_Pad2, CDUXDM, MOUT_n, net_U23032_Pad2, GND, ZOUT_n, net_U23032_Pad2, net_U23030_Pad5, CHWL14_n, WCH14_n, net_U23033_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23034(net_U23030_Pad9, net_U23033_Pad13, net_U23030_Pad8, CH1414, RCH14_n, net_U23030_Pad9, GND, net_U23030_Pad9, F5ASB2_n, CDUYD, XB1_n, net_U23031_Pad12, net_U23032_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23035(CDUYDP, POUT_n, net_U23032_Pad6, CDUYDM, MOUT_n, net_U23032_Pad6, GND, ZOUT_n, net_U23032_Pad6, net_U23030_Pad11, CHWL13_n, WCH14_n, net_U23035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23036(net_U23036_Pad1, net_U23035_Pad13, net_U23036_Pad3, CH1413, RCH14_n, net_U23036_Pad1, GND, net_U23036_Pad1, F5ASB2_n, CDUZD, XB2_n, net_U23031_Pad12, net_U23032_Pad9, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23037(net_U23036_Pad1, CCH14, net_U23037_Pad3, CCH14, net_U23037_Pad5, net_U23037_Pad6, GND, net_U23037_Pad8, net_U23037_Pad9, CCH14, net_U23037_Pad11, net_U23036_Pad3, net_U23037_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23038(CDUZDP, POUT_n, net_U23032_Pad8, CDUZDM, MOUT_n, net_U23032_Pad8, GND, ZOUT_n, net_U23032_Pad8, net_U23037_Pad13, CHWL12_n, WCH14_n, net_U23038_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23039(net_U23037_Pad3, net_U23038_Pad13, net_U23037_Pad6, CH1412, RCH14_n, net_U23037_Pad3, GND, net_U23037_Pad3, F5ASB2_n, TRUND, XB3_n, net_U23031_Pad12, net_U23032_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23040(__A23_2__TRNDP, POUT_n, net_U23032_Pad10, __A23_2__TRNDM, MOUT_n, net_U23032_Pad10, GND, ZOUT_n, net_U23032_Pad10, net_U23037_Pad5, CHWL11_n, WCH14_n, net_U23040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23041(net_U23037_Pad9, net_U23040_Pad13, net_U23037_Pad8, CH1411, RCH14_n, net_U23037_Pad9, GND, net_U23037_Pad9, F5ASB2_n, SHAFTD, XB4_n, net_U23031_Pad12, net_U23032_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23042(__A23_2__SHFTDP, POUT_n, net_U23032_Pad12, __A23_2__SHFTDM, MOUT_n, net_U23032_Pad12, GND, ZOUT_n, net_U23032_Pad12, net_U23037_Pad11, CHWL05_n, __A23_2__WCH07_n, net_U23042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23043(net_U23043_Pad1, net_U23042_Pad13, E5, E5, net_U23043_Pad1, __A23_2__CCH07, GND, __A23_2__RCH07_n, net_U23043_Pad1, CH0705, CHWL06_n, __A23_2__WCH07_n, net_U23043_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23044(net_U23044_Pad1, net_U23043_Pad13, E6, E6, net_U23044_Pad1, __A23_2__CCH07, GND, __A23_2__RCH07_n, net_U23044_Pad1, CH0706, CHWL07_n, __A23_2__WCH07_n, net_U23044_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23045(E7_n, net_U23044_Pad13, net_U23045_Pad3, net_U23045_Pad3, E7_n, __A23_2__CCH07, GND, __A23_2__RCH07_n, E7_n, CH0707, XB7_n, XT0_n, net_U23045_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23046(WCHG_n, XT0_n, CCHG_n, XB7_n, XT0_n, __A23_2__CCH07, GND, net_U23046_Pad8, T6ON_n, T6RPT, CCH13, net_U23046_Pad12, XB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U23047(net_U23046_Pad12, __A23_2__WCH07_n, net_U23045_Pad13, __A23_2__RCH07_n, net_U23047_Pad5, __A23_2__OT1108, GND, __A23_2__OT1113, net_U23047_Pad9, __A23_2__OT1114, net_U23047_Pad11, __A23_2__OT1116, net_U23047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23048(net_U23048_Pad1, CHWL08_n, WCH11_n, net_U23047_Pad5, net_U23048_Pad1, net_U23048_Pad10, GND, net_U23047_Pad5, CCH11, net_U23048_Pad10, RCH11_n, net_U23047_Pad5, CH1108, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23049(net_U23049_Pad1, CHWL13_n, WCH11_n, net_U23047_Pad9, net_U23049_Pad1, net_U23049_Pad10, GND, net_U23047_Pad9, CCH11, net_U23049_Pad10, RCH11_n, net_U23047_Pad9, CH1113, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23050(net_U23050_Pad1, CHWL14_n, WCH11_n, net_U23047_Pad11, net_U23050_Pad1, net_U23050_Pad10, GND, net_U23047_Pad11, CCH11, net_U23050_Pad10, RCH11_n, net_U23047_Pad11, CH1114, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23051(net_U23051_Pad1, CHWL16_n, WCH11_n, net_U23047_Pad13, net_U23051_Pad1, net_U23051_Pad10, GND, net_U23047_Pad13, CCH11, net_U23051_Pad10, RCH11_n, net_U23047_Pad13, CH1116, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23052(net_U23052_Pad1, CHWL16_n, WCH12_n, net_U23052_Pad12, net_U23052_Pad1, net_U23052_Pad10, GND, net_U23052_Pad12, CCH12, net_U23052_Pad10, RCH12_n, net_U23052_Pad12, CH1216, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U23053(net_U23052_Pad12, __A23_2__ISSTDC,  ,  , net_U23053_Pad5, ALTEST, GND, __A23_1__P04A, P04_n, __A23_1__PIPSAM_n, __A23_1__PIPSAM, __A23_1__PIPAXp_n, PIPAXp, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23054(net_U23054_Pad1, CHWL16_n, WCH13_n, T6ON_n, net_U23054_Pad1, net_U23046_Pad8, GND, RCH13_n, T6ON_n, CH1316, CHWL10_n, WCH13_n, net_U23054_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23055(net_U23053_Pad5, net_U23054_Pad13, net_U23055_Pad3, net_U23055_Pad3, net_U23053_Pad5, CCH13, GND, RCH13_n, net_U23053_Pad5, CH1310, __A23_1__PIPSAM_n, __A23_1__PIPAXp_n, __A23_1__PIPGXp, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U23056(PIPAXm, __A23_1__PIPAXm_n, PIPAYp, __A23_1__PIPAYp_n, PIPAYm, __A23_1__PIPAYm_n, GND, __A23_1__PIPAZp_n, PIPAZp, __A23_1__PIPAZm_n, PIPAZm,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23057(__A23_1__PIPGXm, __A23_1__PIPSAM_n, __A23_1__PIPAXm_n, __A23_1__PIPGYp, __A23_1__PIPSAM_n, __A23_1__PIPAYp_n, GND, __A23_1__PIPSAM_n, __A23_1__PIPAYm_n, __A23_1__PIPGYm, __A23_1__PIPSAM_n, __A23_1__PIPAZp_n, __A23_1__PIPGZp, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23058(__A23_1__PIPGZm, __A23_1__PIPSAM_n, __A23_1__PIPAZm_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule