`timescale 1ns/1ps
`default_nettype none

module four_bit_1(SIM_RST, SIM_CLK, p4VSW, GND, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI01_n, MONEX, PONEX, TWOX, XUY05_n, XUY06_n, CH01, CH02, CH03, CH04, G01ED, G02ED, G03ED, G04ED, MCRO_n, G2LSG_n, G05_n, G06_n, G07_n, MDT01, MDT02, MDT03, MDT04, SA01, SA02, SA03, SA04, RBLG_n, RULOG_n, WL05_n, WL06_n, WG1G_n, WG3G_n, WG4G_n, WYDLOG_n, WYDG_n, WYLOG_n, RB1, R1C, R15, RB2, WL16_n, WHOMP, WHOMPA, CI05_n, CO06, G01, G01_n, G02, G03, G04, L01_n, L02_n, L04_n, RL01_n, RL02_n, RL03_n, RL04_n, SUMA01_n, SUMB01_n, SUMA02_n, SUMB02_n, SUMA03_n, SUMB03_n, WL01, WL01_n, WL02, WL02_n, WL03, WL03_n, WL04, WL04_n, XUY01_n, XUY02_n, GEM01, GEM02, GEM03, GEM04, MWL01, MWL02, MWL03, MWL04);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire A2XG_n;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH01;
    input wire CH02;
    input wire CH03;
    input wire CH04;
    input wire CI01_n;
    output wire CI05_n;
    input wire CLG1G;
    input wire CLXC;
    output wire CO06; //FPGA#wand
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire G01;
    input wire G01ED;
    inout wire G01_n; //FPGA#wand
    output wire G02;
    input wire G02ED;
    output wire G03;
    input wire G03ED;
    output wire G04;
    input wire G04ED;
    input wire G05_n;
    input wire G06_n;
    input wire G07_n;
    input wire G2LSG_n;
    output wire GEM01;
    output wire GEM02;
    output wire GEM03;
    output wire GEM04;
    inout wire L01_n; //FPGA#wand
    inout wire L02_n; //FPGA#wand
    inout wire L04_n; //FPGA#wand
    input wire L2GDG_n;
    input wire MCRO_n;
    input wire MDT01;
    input wire MDT02;
    input wire MDT03;
    input wire MDT04;
    input wire MONEX;
    output wire MWL01; //FPGA#wand
    output wire MWL02; //FPGA#wand
    output wire MWL03; //FPGA#wand
    output wire MWL04; //FPGA#wand
    input wire PONEX;
    input wire R15;
    input wire R1C;
    input wire RAG_n;
    input wire RB1;
    input wire RB2;
    input wire RBLG_n;
    input wire RCG_n;
    input wire RGG_n;
    inout wire RL01_n; //FPGA#wand
    inout wire RL02_n; //FPGA#wand
    inout wire RL03_n; //FPGA#wand
    inout wire RL04_n; //FPGA#wand
    input wire RLG_n;
    input wire RQG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA01;
    input wire SA02;
    input wire SA03;
    input wire SA04;
    output wire SUMA01_n;
    output wire SUMA02_n;
    output wire SUMA03_n;
    output wire SUMB01_n;
    output wire SUMB02_n;
    output wire SUMB03_n;
    input wire TWOX;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WHOMP;
    input wire WHOMPA;
    output wire WL01;
    output wire WL01_n;
    output wire WL02;
    output wire WL02_n;
    output wire WL03;
    output wire WL03_n;
    output wire WL04;
    output wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL16_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYDLOG_n;
    input wire WYLOG_n;
    input wire WZG_n;
    output wire XUY01_n;
    output wire XUY02_n;
    input wire XUY05_n;
    input wire XUY06_n;
    wire __A08_1__X1;
    wire __A08_1__X1_n;
    wire __A08_1__X2;
    wire __A08_1__X2_n;
    wire __A08_1__Y1;
    wire __A08_1__Y1_n;
    wire __A08_1__Y2;
    wire __A08_1__Y2_n;
    wire __A08_1___A1_n;
    wire __A08_1___A2_n;
    wire __A08_1___B1_n;
    wire __A08_1___B2_n;
    wire __A08_1___CI_INTERNAL;
    wire __A08_1___G2_n; //FPGA#wand
    wire __A08_1___Q1_n;
    wire __A08_1___Q2_n;
    wire __A08_1___RL_OUT_1;
    wire __A08_1___RL_OUT_2;
    wire __A08_1___Z1_n; //FPGA#wand
    wire __A08_1___Z2_n; //FPGA#wand
    wire __A08_2__X1;
    wire __A08_2__X1_n;
    wire __A08_2__X2;
    wire __A08_2__X2_n;
    wire __A08_2__Y1;
    wire __A08_2__Y1_n;
    wire __A08_2__Y2;
    wire __A08_2__Y2_n;
    wire __A08_2___A1_n;
    wire __A08_2___A2_n;
    wire __A08_2___B1_n;
    wire __A08_2___B2_n;
    wire __A08_2___CI_INTERNAL;
    wire __A08_2___G1_n; //FPGA#wand
    wire __A08_2___Q1_n;
    wire __A08_2___Q2_n;
    wire __A08_2___RL_OUT_1;
    wire __A08_2___RL_OUT_2;
    wire __A08_2___SUMA2;
    wire __A08_2___SUMB2;
    wire __A08_2___Z1_n; //FPGA#wand
    wire __A08_2___Z2_n; //FPGA#wand
    wire __CI03_n;
    wire __CO04; //FPGA#wand
    wire __G04_n; //FPGA#wand
    wire __L03_n; //FPGA#wand
    wire __XUY03_n;
    wire __XUY04_n;
    wire net_U8001_Pad1;
    wire net_U8001_Pad10;
    wire net_U8001_Pad4;
    wire net_U8003_Pad1;
    wire net_U8003_Pad10;
    wire net_U8004_Pad1;
    wire net_U8004_Pad12;
    wire net_U8004_Pad13;
    wire net_U8004_Pad2;
    wire net_U8004_Pad6;
    wire net_U8004_Pad8;
    wire net_U8005_Pad12;
    wire net_U8005_Pad2;
    wire net_U8006_Pad10;
    wire net_U8006_Pad13;
    wire net_U8006_Pad4;
    wire net_U8007_Pad11;
    wire net_U8007_Pad13;
    wire net_U8007_Pad3;
    wire net_U8007_Pad5;
    wire net_U8007_Pad9;
    wire net_U8008_Pad1;
    wire net_U8008_Pad10;
    wire net_U8008_Pad13;
    wire net_U8008_Pad4;
    wire net_U8009_Pad1;
    wire net_U8009_Pad13;
    wire net_U8009_Pad4;
    wire net_U8010_Pad1;
    wire net_U8010_Pad13;
    wire net_U8010_Pad4;
    wire net_U8011_Pad10;
    wire net_U8011_Pad11;
    wire net_U8011_Pad13;
    wire net_U8011_Pad8;
    wire net_U8011_Pad9;
    wire net_U8012_Pad13;
    wire net_U8012_Pad4;
    wire net_U8013_Pad1;
    wire net_U8013_Pad11;
    wire net_U8013_Pad13;
    wire net_U8013_Pad5;
    wire net_U8013_Pad9;
    wire net_U8014_Pad10;
    wire net_U8014_Pad13;
    wire net_U8016_Pad1;
    wire net_U8016_Pad4;
    wire net_U8018_Pad11;
    wire net_U8018_Pad12;
    wire net_U8018_Pad13;
    wire net_U8019_Pad1;
    wire net_U8019_Pad10;
    wire net_U8019_Pad4;
    wire net_U8021_Pad1;
    wire net_U8021_Pad13;
    wire net_U8022_Pad1;
    wire net_U8022_Pad12;
    wire net_U8022_Pad8;
    wire net_U8023_Pad10;
    wire net_U8023_Pad13;
    wire net_U8023_Pad4;
    wire net_U8024_Pad10;
    wire net_U8024_Pad11;
    wire net_U8024_Pad4;
    wire net_U8024_Pad9;
    wire net_U8026_Pad4;
    wire net_U8026_Pad5;
    wire net_U8026_Pad6;
    wire net_U8026_Pad8;
    wire net_U8027_Pad1;
    wire net_U8027_Pad10;
    wire net_U8028_Pad13;
    wire net_U8028_Pad3;
    wire net_U8028_Pad9;
    wire net_U8029_Pad1;
    wire net_U8029_Pad10;
    wire net_U8030_Pad1;
    wire net_U8030_Pad10;
    wire net_U8030_Pad13;
    wire net_U8031_Pad13;
    wire net_U8031_Pad2;
    wire net_U8031_Pad3;
    wire net_U8031_Pad4;
    wire net_U8031_Pad8;
    wire net_U8035_Pad1;
    wire net_U8035_Pad10;
    wire net_U8035_Pad4;
    wire net_U8037_Pad1;
    wire net_U8037_Pad10;
    wire net_U8038_Pad1;
    wire net_U8038_Pad12;
    wire net_U8038_Pad2;
    wire net_U8038_Pad6;
    wire net_U8038_Pad8;
    wire net_U8039_Pad12;
    wire net_U8039_Pad2;
    wire net_U8040_Pad10;
    wire net_U8040_Pad13;
    wire net_U8040_Pad4;
    wire net_U8041_Pad11;
    wire net_U8041_Pad13;
    wire net_U8041_Pad3;
    wire net_U8041_Pad5;
    wire net_U8041_Pad9;
    wire net_U8042_Pad10;
    wire net_U8042_Pad11;
    wire net_U8042_Pad4;
    wire net_U8042_Pad9;
    wire net_U8044_Pad1;
    wire net_U8044_Pad6;
    wire net_U8045_Pad13;
    wire net_U8045_Pad4;
    wire net_U8046_Pad1;
    wire net_U8046_Pad13;
    wire net_U8046_Pad4;
    wire net_U8047_Pad1;
    wire net_U8047_Pad13;
    wire net_U8047_Pad4;
    wire net_U8048_Pad1;
    wire net_U8048_Pad10;
    wire net_U8048_Pad13;
    wire net_U8048_Pad4;
    wire net_U8049_Pad11;
    wire net_U8049_Pad8;
    wire net_U8050_Pad11;
    wire net_U8050_Pad13;
    wire net_U8050_Pad5;
    wire net_U8052_Pad11;
    wire net_U8052_Pad12;
    wire net_U8052_Pad13;
    wire net_U8053_Pad1;
    wire net_U8053_Pad10;
    wire net_U8053_Pad4;
    wire net_U8055_Pad13;
    wire net_U8056_Pad10;
    wire net_U8056_Pad13;
    wire net_U8056_Pad4;
    wire net_U8057_Pad10;
    wire net_U8057_Pad11;
    wire net_U8057_Pad4;
    wire net_U8057_Pad9;
    wire net_U8059_Pad4;
    wire net_U8059_Pad5;
    wire net_U8059_Pad6;
    wire net_U8059_Pad8;
    wire net_U8060_Pad1;
    wire net_U8060_Pad10;
    wire net_U8061_Pad3;
    wire net_U8062_Pad1;
    wire net_U8062_Pad10;
    wire net_U8063_Pad1;
    wire net_U8063_Pad10;

    pullup R8001(__CO04);
    pullup R8002(RL01_n);
    pullup R8003(L01_n);
    pullup R8005(__A08_1___Z1_n);
    pullup R8006(G01_n);
    pullup R8007(RL02_n);
    pullup R8008(L02_n);
    pullup R8009(__A08_1___Z2_n);
    pullup R8010(__A08_1___G2_n);
    pullup R8011(CO06);
    pullup R8012(RL03_n);
    pullup R8013(__L03_n);
    pullup R8015(__A08_2___Z1_n);
    pullup R8016(__A08_2___G1_n);
    pullup R8017(RL04_n);
    pullup R8018(L04_n);
    pullup R8019(__A08_2___Z2_n);
    pullup R8020(__G04_n);
    U74HC02 U8001(net_U8001_Pad1, A2XG_n, __A08_1___A1_n, net_U8001_Pad4, WYLOG_n, WL01_n, GND, WL16_n, WYDLOG_n, net_U8001_Pad10, __A08_1__Y1_n, CUG, __A08_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8002(PONEX, net_U8001_Pad1, __A08_1__X1_n, CLXC, CUG, __A08_1__X1, GND, __A08_1__Y1_n, net_U8001_Pad4, net_U8001_Pad10, __A08_1__Y1, __A08_1__X1_n, __A08_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8003(net_U8003_Pad1, __A08_1__X1_n, __A08_1__Y1_n, XUY01_n, __A08_1__X1, __A08_1__Y1, GND, net_U8003_Pad1, XUY01_n, net_U8003_Pad10, net_U8003_Pad1, SUMA01_n, __A08_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8004(net_U8004_Pad1, net_U8004_Pad2, SUMA01_n, SUMB01_n, RULOG_n, net_U8004_Pad6, GND, net_U8004_Pad8, __XUY03_n, XUY01_n, CI01_n, net_U8004_Pad12, net_U8004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8005(CI01_n, net_U8005_Pad2, G01_n, GEM01, RL01_n, WL01, GND, WL01_n, WL01,  ,  , net_U8005_Pad12, __A08_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8006(SUMB01_n, net_U8003_Pad10, net_U8005_Pad2, net_U8006_Pad4, WAG_n, WL01_n, GND, WL03_n, WALSG_n, net_U8006_Pad10, __A08_1___A1_n, CAG, net_U8006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8007(net_U8004_Pad8, __CO04, net_U8007_Pad3, RL01_n, net_U8007_Pad5, L01_n, GND, __A08_1___Z1_n, net_U8007_Pad9, RL01_n, net_U8007_Pad11, RL01_n, net_U8007_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U8008(net_U8008_Pad1, RAG_n, __A08_1___A1_n, net_U8008_Pad4, WLG_n, WL01_n, GND, __G04_n, G2LSG_n, net_U8008_Pad10, L01_n, CLG1G, net_U8008_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8009(net_U8009_Pad1, WG1G_n, WL04_n, net_U8009_Pad4, WQG_n, WL01_n, GND, net_U8009_Pad4, net_U8009_Pad13, __A08_1___Q1_n, __A08_1___Q1_n, CQG, net_U8009_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8010(net_U8010_Pad1, RQG_n, __A08_1___Q1_n, net_U8010_Pad4, WZG_n, WL01_n, GND, net_U8010_Pad4, net_U8010_Pad13, net_U8007_Pad9, __A08_1___Z1_n, CZG, net_U8010_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8011(__A08_1___RL_OUT_1, net_U8010_Pad1, MDT01, RB1, R15, net_U8007_Pad13, GND, net_U8011_Pad8, net_U8011_Pad9, net_U8011_Pad10, net_U8011_Pad11, net_U8007_Pad11, net_U8011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8012(net_U8011_Pad13, RZG_n, __A08_1___Z1_n, net_U8012_Pad4, WBG_n, WL01_n, GND, net_U8012_Pad4, net_U8012_Pad13, __A08_1___B1_n, __A08_1___B1_n, CBG, net_U8012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8013(net_U8013_Pad1, __CO04, net_U8011_Pad8, RL01_n, net_U8013_Pad5, G01_n, GND, G01_n, net_U8013_Pad9, RL02_n, net_U8013_Pad11, L02_n, net_U8013_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U8014(net_U8011_Pad9, RBLG_n, __A08_1___B1_n, net_U8011_Pad10, net_U8012_Pad13, RCG_n, GND, WL16_n, WG3G_n, net_U8014_Pad10, WL02_n, WG4G_n, net_U8014_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8015(net_U8006_Pad4, net_U8006_Pad10, net_U8004_Pad6, net_U8008_Pad1, CH01, net_U8007_Pad3, GND, net_U8007_Pad5, net_U8008_Pad4, net_U8008_Pad10, net_U8008_Pad13, __A08_1___A1_n, net_U8006_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8016(net_U8016_Pad1, L2GDG_n, MCRO_n, net_U8016_Pad4, WG1G_n, WL01_n, GND, G01_n, CGG, G01, RGG_n, G01_n, net_U8011_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8017(net_U8016_Pad1, net_U8016_Pad4, WHOMPA, __XUY04_n, XUY02_n, net_U8013_Pad1, GND, __A08_1___RL_OUT_1, RLG_n, L01_n, GND, net_U8013_Pad9, G01, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U8018(net_U8013_Pad5, G01ED, SA01, net_U8014_Pad10, net_U8014_Pad13,  , GND,  , G02ED, SA02, net_U8018_Pad11, net_U8018_Pad12, net_U8018_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8019(net_U8019_Pad1, A2XG_n, __A08_1___A2_n, net_U8019_Pad4, WYLOG_n, WL02_n, GND, WL01_n, WYDG_n, net_U8019_Pad10, __A08_1__Y2_n, CUG, __A08_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8020(TWOX, net_U8019_Pad1, __A08_1__X2_n, CLXC, CUG, __A08_1__X2, GND, __A08_1__Y2_n, net_U8019_Pad4, net_U8019_Pad10, __A08_1__Y2, __A08_1__X2_n, __A08_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8021(net_U8021_Pad1, __A08_1__X2_n, __A08_1__Y2_n, XUY02_n, __A08_1__X2, __A08_1__Y2, GND, __G04_n, CGG, G04, net_U8021_Pad1, XUY02_n, net_U8021_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8022(net_U8022_Pad1, net_U8009_Pad1, net_U8021_Pad1, SUMA02_n, GND, __CI03_n, GND, net_U8022_Pad8, SUMA02_n, SUMB02_n, RULOG_n, net_U8022_Pad12, G04, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8023(SUMB02_n, net_U8021_Pad13, net_U8005_Pad12, net_U8023_Pad4, WAG_n, WL02_n, GND, WL04_n, WALSG_n, net_U8023_Pad10, __A08_1___A2_n, CAG, net_U8023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8024(net_U8023_Pad4, net_U8023_Pad10, net_U8022_Pad8, net_U8024_Pad4, CH02, net_U8013_Pad11, GND, net_U8013_Pad13, net_U8024_Pad9, net_U8024_Pad10, net_U8024_Pad11, __A08_1___A2_n, net_U8023_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8025(net_U8024_Pad4, RAG_n, __A08_1___A2_n, net_U8024_Pad9, WLG_n, WL02_n, GND, G05_n, G2LSG_n, net_U8024_Pad10, L02_n, CLG1G, net_U8024_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8026(RLG_n, L02_n, __A08_1___RL_OUT_2, net_U8026_Pad4, net_U8026_Pad5, net_U8026_Pad6, GND, net_U8026_Pad8, MDT02, R1C, RB2, __A08_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8027(net_U8027_Pad1, WQG_n, WL02_n, __A08_1___Q2_n, net_U8027_Pad1, net_U8027_Pad10, GND, __A08_1___Q2_n, CQG, net_U8027_Pad10, RQG_n, __A08_1___Q2_n, net_U8026_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8028(net_U8026_Pad6, RL02_n, net_U8028_Pad3, __A08_1___Z2_n, net_U8026_Pad8, RL02_n, GND, RL02_n, net_U8028_Pad9, __A08_1___G2_n, net_U8018_Pad13, __A08_1___G2_n, net_U8028_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8029(net_U8029_Pad1, WZG_n, WL02_n, net_U8028_Pad3, net_U8029_Pad1, net_U8029_Pad10, GND, __A08_1___Z2_n, CZG, net_U8029_Pad10, RZG_n, __A08_1___Z2_n, net_U8026_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8030(net_U8030_Pad1, WBG_n, WL02_n, __A08_1___B2_n, net_U8030_Pad1, net_U8030_Pad10, GND, __A08_1___B2_n, CBG, net_U8030_Pad10, RBLG_n, __A08_1___B2_n, net_U8030_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U8031(net_U8030_Pad13, net_U8031_Pad2, net_U8031_Pad3, net_U8031_Pad4, G02, net_U8028_Pad13, GND, net_U8031_Pad8, GND, XUY06_n, __XUY04_n, net_U8028_Pad9, net_U8031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8032(net_U8031_Pad2, net_U8030_Pad10, RCG_n, net_U8018_Pad11, WL01_n, WG3G_n, GND, WL03_n, WG4G_n, net_U8018_Pad12, L2GDG_n, L01_n, net_U8031_Pad3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8033(net_U8031_Pad4, WG1G_n, WL02_n, G02, __A08_1___G2_n, CGG, GND, RGG_n, __A08_1___G2_n, net_U8031_Pad13, RGG_n, __G04_n, net_U8004_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8034(__A08_1___G2_n, GEM02, RL02_n, WL02, WL02, WL02_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8035(net_U8035_Pad1, A2XG_n, __A08_2___A1_n, net_U8035_Pad4, WYLOG_n, WL03_n, GND, WL02_n, WYDG_n, net_U8035_Pad10, __A08_2__Y1_n, CUG, __A08_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8036(MONEX, net_U8035_Pad1, __A08_2__X1_n, CLXC, CUG, __A08_2__X1, GND, __A08_2__Y1_n, net_U8035_Pad4, net_U8035_Pad10, __A08_2__Y1, __A08_2__X1_n, __A08_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8037(net_U8037_Pad1, __A08_2__X1_n, __A08_2__Y1_n, __XUY03_n, __A08_2__X1, __A08_2__Y1, GND, net_U8037_Pad1, __XUY03_n, net_U8037_Pad10, net_U8037_Pad1, SUMA03_n, __A08_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8038(net_U8038_Pad1, net_U8038_Pad2, SUMA03_n, SUMB03_n, RULOG_n, net_U8038_Pad6, GND, net_U8038_Pad8, XUY05_n, __XUY03_n, __CI03_n, net_U8038_Pad12, G03, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8039(__CI03_n, net_U8039_Pad2, __A08_2___G1_n, GEM03, RL03_n, WL03, GND, WL03_n, WL03,  ,  , net_U8039_Pad12, __A08_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8040(SUMB03_n, net_U8037_Pad10, net_U8039_Pad2, net_U8040_Pad4, WAG_n, WL03_n, GND, WL05_n, WALSG_n, net_U8040_Pad10, __A08_2___A1_n, CAG, net_U8040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8041(net_U8038_Pad8, CO06, net_U8041_Pad3, RL03_n, net_U8041_Pad5, __L03_n, GND, __A08_2___Z1_n, net_U8041_Pad9, RL03_n, net_U8041_Pad11, RL03_n, net_U8041_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1) U8042(net_U8040_Pad4, net_U8040_Pad10, net_U8038_Pad6, net_U8042_Pad4, CH03, net_U8041_Pad3, GND, net_U8041_Pad5, net_U8042_Pad9, net_U8042_Pad10, net_U8042_Pad11, __A08_2___A1_n, net_U8040_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8043(net_U8042_Pad4, RAG_n, __A08_2___A1_n, net_U8042_Pad9, WLG_n, WL03_n, GND, G06_n, G2LSG_n, net_U8042_Pad10, __L03_n, CLG1G, net_U8042_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8044(net_U8044_Pad1, __A08_2___SUMA2, __A08_2___SUMA2, __A08_2___SUMB2, RULOG_n, net_U8044_Pad6, GND, __A08_2___RL_OUT_1, RLG_n, __L03_n, GND, CI05_n, __CO04, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8045( ,  ,  , net_U8045_Pad4, WQG_n, WL03_n, GND, net_U8045_Pad4, net_U8045_Pad13, __A08_2___Q1_n, __A08_2___Q1_n, CQG, net_U8045_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8046(net_U8046_Pad1, RQG_n, __A08_2___Q1_n, net_U8046_Pad4, WZG_n, WL03_n, GND, net_U8046_Pad4, net_U8046_Pad13, net_U8041_Pad9, __A08_2___Z1_n, CZG, net_U8046_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8047(net_U8047_Pad1, RZG_n, __A08_2___Z1_n, net_U8047_Pad4, WBG_n, WL03_n, GND, net_U8047_Pad4, net_U8047_Pad13, __A08_2___B1_n, __A08_2___B1_n, CBG, net_U8047_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8048(net_U8048_Pad1, RBLG_n, __A08_2___B1_n, net_U8048_Pad4, net_U8047_Pad13, RCG_n, GND, WL02_n, WG3G_n, net_U8048_Pad10, WL04_n, WG4G_n, net_U8048_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8049(__A08_2___RL_OUT_1, net_U8046_Pad1, MDT03, R1C, R15, net_U8041_Pad13, GND, net_U8049_Pad8, net_U8048_Pad1, net_U8048_Pad4, net_U8049_Pad11, net_U8041_Pad11, net_U8047_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8050(net_U8031_Pad8, CO06, net_U8049_Pad8, RL03_n, net_U8050_Pad5, __A08_2___G1_n, GND, __A08_2___G1_n, net_U8038_Pad12, RL04_n, net_U8050_Pad11, L04_n, net_U8050_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U8051(net_U8038_Pad1, L2GDG_n, L02_n, net_U8038_Pad2, WG1G_n, WL03_n, GND, __A08_2___G1_n, CGG, G03, RGG_n, __A08_2___G1_n, net_U8049_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U8052(net_U8050_Pad5, G03ED, SA03, net_U8048_Pad10, net_U8048_Pad13,  , GND,  , G04ED, SA04, net_U8052_Pad11, net_U8052_Pad12, net_U8052_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8053(net_U8053_Pad1, A2XG_n, __A08_2___A2_n, net_U8053_Pad4, WYLOG_n, WL04_n, GND, WL03_n, WYDG_n, net_U8053_Pad10, __A08_2__Y2_n, CUG, __A08_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8054(MONEX, net_U8053_Pad1, __A08_2__X2_n, CLXC, CUG, __A08_2__X2, GND, __A08_2__Y2_n, net_U8053_Pad4, net_U8053_Pad10, __A08_2__Y2, __A08_2__X2_n, __A08_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8055(net_U8044_Pad1, __A08_2__X2_n, __A08_2__Y2_n, __XUY04_n, __A08_2__X2, __A08_2__Y2, GND,  ,  ,  , net_U8044_Pad1, __XUY04_n, net_U8055_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8056(__A08_2___SUMB2, net_U8055_Pad13, net_U8039_Pad12, net_U8056_Pad4, WAG_n, WL04_n, GND, WL06_n, WALSG_n, net_U8056_Pad10, __A08_2___A2_n, CAG, net_U8056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8057(net_U8056_Pad4, net_U8056_Pad10, net_U8044_Pad6, net_U8057_Pad4, CH04, net_U8050_Pad11, GND, net_U8050_Pad13, net_U8057_Pad9, net_U8057_Pad10, net_U8057_Pad11, __A08_2___A2_n, net_U8056_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8058(net_U8057_Pad4, RAG_n, __A08_2___A2_n, net_U8057_Pad9, WLG_n, WL04_n, GND, G07_n, G2LSG_n, net_U8057_Pad10, L04_n, CLG1G, net_U8057_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8059(RLG_n, L04_n, __A08_2___RL_OUT_2, net_U8059_Pad4, net_U8059_Pad5, net_U8059_Pad6, GND, net_U8059_Pad8, MDT04, R1C, R15, __A08_2___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8060(net_U8060_Pad1, WQG_n, WL04_n, __A08_2___Q2_n, net_U8060_Pad1, net_U8060_Pad10, GND, __A08_2___Q2_n, CQG, net_U8060_Pad10, RQG_n, __A08_2___Q2_n, net_U8059_Pad4, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8061(net_U8059_Pad6, RL04_n, net_U8061_Pad3, __A08_2___Z2_n, net_U8059_Pad8, RL04_n, GND, RL04_n, net_U8004_Pad12, __G04_n, net_U8052_Pad13, __G04_n, net_U8022_Pad12, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8062(net_U8062_Pad1, WZG_n, WL04_n, net_U8061_Pad3, net_U8062_Pad1, net_U8062_Pad10, GND, __A08_2___Z2_n, CZG, net_U8062_Pad10, RZG_n, __A08_2___Z2_n, net_U8059_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8063(net_U8063_Pad1, WBG_n, WL04_n, __A08_2___B2_n, net_U8063_Pad1, net_U8063_Pad10, GND, __A08_2___B2_n, CBG, net_U8063_Pad10, RBLG_n, __A08_2___B2_n, net_U8004_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8064(net_U8004_Pad2, net_U8063_Pad10, RCG_n, net_U8052_Pad11, WL03_n, WG3G_n, GND, WL05_n, WG4G_n, net_U8052_Pad12, L2GDG_n, __L03_n, net_U8022_Pad1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8065(__G04_n, GEM04, RL04_n, WL04, WL04, WL04_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U8066(SUMA01_n, net_U8003_Pad1, XUY01_n, CI01_n, GND,  , GND,  , net_U8021_Pad1, XUY02_n, __A08_1___CI_INTERNAL, WHOMP, SUMA02_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U8067(SUMA03_n, net_U8037_Pad1, __XUY03_n, __CI03_n, GND,  , GND,  , net_U8044_Pad1, __XUY04_n, __A08_2___CI_INTERNAL, WHOMP, __A08_2___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U8068(RL01_n, MWL01, RL02_n, MWL02, RL03_n, MWL03, GND, MWL04, RL04_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8
endmodule